<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-57.3194,161.541,175.044,41.7</PageViewport>
<gate>
<ID>193</ID>
<type>AE_SMALL_INVERTER</type>
<position>69,110</position>
<input>
<ID>IN_0</ID>92 </input>
<output>
<ID>OUT_0</ID>97 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>194</ID>
<type>AE_SMALL_INVERTER</type>
<position>69,118</position>
<input>
<ID>IN_0</ID>93 </input>
<output>
<ID>OUT_0</ID>96 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>195</ID>
<type>AE_SMALL_INVERTER</type>
<position>69,126</position>
<input>
<ID>IN_0</ID>94 </input>
<output>
<ID>OUT_0</ID>98 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>196</ID>
<type>AE_SMALL_INVERTER</type>
<position>69,134</position>
<input>
<ID>IN_0</ID>95 </input>
<output>
<ID>OUT_0</ID>99 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>197</ID>
<type>AA_TOGGLE</type>
<position>92,64</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>198</ID>
<type>AA_LABEL</type>
<position>92,61.5</position>
<gparam>LABEL_TEXT S3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>AA_TOGGLE</type>
<position>71,143</position>
<output>
<ID>OUT_0</ID>95 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_TOGGLE</type>
<position>74,143</position>
<output>
<ID>OUT_0</ID>94 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>406</ID>
<type>AA_LABEL</type>
<position>57,160</position>
<gparam>LABEL_TEXT Unidade Aritmetica</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>AA_TOGGLE</type>
<position>77,143</position>
<output>
<ID>OUT_0</ID>93 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_TOGGLE</type>
<position>80,143</position>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>410</ID>
<type>AA_LABEL</type>
<position>61,141</position>
<gparam>LABEL_TEXT 74HC08</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>411</ID>
<type>AA_LABEL</type>
<position>52.5,139</position>
<gparam>LABEL_TEXT 74HC32</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>AA_TOGGLE</type>
<position>83,143</position>
<output>
<ID>OUT_0</ID>91 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>412</ID>
<type>AA_LABEL</type>
<position>69.5,75</position>
<gparam>LABEL_TEXT 74HC04</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>413</ID>
<type>AA_LABEL</type>
<position>52.5,132</position>
<gparam>LABEL_TEXT U1a</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>AA_TOGGLE</type>
<position>86,143</position>
<output>
<ID>OUT_0</ID>89 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>414</ID>
<type>AA_LABEL</type>
<position>52.5,124</position>
<gparam>LABEL_TEXT U1b</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>415</ID>
<type>AA_LABEL</type>
<position>52.5,116</position>
<gparam>LABEL_TEXT U1c</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>AA_TOGGLE</type>
<position>89,143</position>
<output>
<ID>OUT_0</ID>87 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>416</ID>
<type>AA_LABEL</type>
<position>52.5,108</position>
<gparam>LABEL_TEXT U1d</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>417</ID>
<type>AA_LABEL</type>
<position>52.5,100</position>
<gparam>LABEL_TEXT U1e</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>AA_TOGGLE</type>
<position>92,143</position>
<output>
<ID>OUT_0</ID>83 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>418</ID>
<type>AA_LABEL</type>
<position>52.5,92</position>
<gparam>LABEL_TEXT U1f</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>419</ID>
<type>AA_LABEL</type>
<position>52.5,84</position>
<gparam>LABEL_TEXT U1g</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AA_LABEL</type>
<position>17,145.5</position>
<gparam>LABEL_TEXT X7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>420</ID>
<type>AA_LABEL</type>
<position>52.5,76</position>
<gparam>LABEL_TEXT U1h</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>AA_LABEL</type>
<position>20,145.5</position>
<gparam>LABEL_TEXT X6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>AA_LABEL</type>
<position>23,145.5</position>
<gparam>LABEL_TEXT X5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>422</ID>
<type>AA_LABEL</type>
<position>65.5,137</position>
<gparam>LABEL_TEXT U2a</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>37</ID>
<type>AA_LABEL</type>
<position>26,145.5</position>
<gparam>LABEL_TEXT X4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>423</ID>
<type>AA_LABEL</type>
<position>65.5,133</position>
<gparam>LABEL_TEXT U2b</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>AA_LABEL</type>
<position>29,145.5</position>
<gparam>LABEL_TEXT X3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>424</ID>
<type>AA_LABEL</type>
<position>65.5,129</position>
<gparam>LABEL_TEXT U2c</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>AA_LABEL</type>
<position>32,145.5</position>
<gparam>LABEL_TEXT X2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>425</ID>
<type>AA_LABEL</type>
<position>65.5,125</position>
<gparam>LABEL_TEXT U2d</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>AA_LABEL</type>
<position>35,145.5</position>
<gparam>LABEL_TEXT X1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>426</ID>
<type>AA_LABEL</type>
<position>65.5,121</position>
<gparam>LABEL_TEXT U2e</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>41</ID>
<type>AA_LABEL</type>
<position>38,145.5</position>
<gparam>LABEL_TEXT X0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>427</ID>
<type>AA_LABEL</type>
<position>65.5,117</position>
<gparam>LABEL_TEXT U2f</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>AA_LABEL</type>
<position>71,145.5</position>
<gparam>LABEL_TEXT Y7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>428</ID>
<type>AA_LABEL</type>
<position>65.5,113</position>
<gparam>LABEL_TEXT U2g</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>43</ID>
<type>AA_LABEL</type>
<position>74,145.5</position>
<gparam>LABEL_TEXT Y6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>429</ID>
<type>AA_LABEL</type>
<position>65.5,109</position>
<gparam>LABEL_TEXT U2h</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>44</ID>
<type>AA_LABEL</type>
<position>77,145.5</position>
<gparam>LABEL_TEXT Y5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>430</ID>
<type>AA_LABEL</type>
<position>65.5,105</position>
<gparam>LABEL_TEXT U2i</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>AA_LABEL</type>
<position>80,145.5</position>
<gparam>LABEL_TEXT Y4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>431</ID>
<type>AA_LABEL</type>
<position>65.5,101</position>
<gparam>LABEL_TEXT U2j</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>46</ID>
<type>AA_LABEL</type>
<position>83,145.5</position>
<gparam>LABEL_TEXT Y3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>432</ID>
<type>AA_LABEL</type>
<position>65.5,97</position>
<gparam>LABEL_TEXT U2k</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>47</ID>
<type>AA_LABEL</type>
<position>86,145.5</position>
<gparam>LABEL_TEXT Y2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>433</ID>
<type>AA_LABEL</type>
<position>65.5,93</position>
<gparam>LABEL_TEXT U2l</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>AA_LABEL</type>
<position>89,145.5</position>
<gparam>LABEL_TEXT Y1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>434</ID>
<type>AA_LABEL</type>
<position>65.5,89</position>
<gparam>LABEL_TEXT U2m</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>49</ID>
<type>AA_LABEL</type>
<position>92,145.5</position>
<gparam>LABEL_TEXT Y0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>435</ID>
<type>AA_LABEL</type>
<position>65.5,85</position>
<gparam>LABEL_TEXT U2n</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>436</ID>
<type>AA_LABEL</type>
<position>65.5,81</position>
<gparam>LABEL_TEXT U2o</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>437</ID>
<type>AA_LABEL</type>
<position>65.5,77</position>
<gparam>LABEL_TEXT U2p</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>438</ID>
<type>AA_LABEL</type>
<position>72.5,134</position>
<gparam>LABEL_TEXT U3a</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>439</ID>
<type>AA_LABEL</type>
<position>72.5,126</position>
<gparam>LABEL_TEXT U3b</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>440</ID>
<type>AA_LABEL</type>
<position>72.5,118</position>
<gparam>LABEL_TEXT U3c</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>441</ID>
<type>AA_LABEL</type>
<position>72.5,110</position>
<gparam>LABEL_TEXT U3d</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>442</ID>
<type>AA_LABEL</type>
<position>72.5,102</position>
<gparam>LABEL_TEXT U3e</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>443</ID>
<type>AA_LABEL</type>
<position>72.5,94</position>
<gparam>LABEL_TEXT U3f</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>58</ID>
<type>AA_LABEL</type>
<position>32.5,46.5</position>
<gparam>LABEL_TEXT G3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>444</ID>
<type>AA_LABEL</type>
<position>72.5,86</position>
<gparam>LABEL_TEXT U3g</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>59</ID>
<type>AA_LABEL</type>
<position>35.5,46.5</position>
<gparam>LABEL_TEXT G2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>445</ID>
<type>AA_LABEL</type>
<position>72.5,78</position>
<gparam>LABEL_TEXT U3h</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>AA_LABEL</type>
<position>38.5,46.5</position>
<gparam>LABEL_TEXT G1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>446</ID>
<type>AA_LABEL</type>
<position>27.5,149</position>
<gparam>LABEL_TEXT Entradas (X)</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>61</ID>
<type>AA_LABEL</type>
<position>41.5,46.5</position>
<gparam>LABEL_TEXT G0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>448</ID>
<type>AA_LABEL</type>
<position>81.5,149</position>
<gparam>LABEL_TEXT Entradas (Y)</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>449</ID>
<type>AA_LABEL</type>
<position>28.5,43.5</position>
<gparam>LABEL_TEXT Saidas (G)</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>450</ID>
<type>AA_LABEL</type>
<position>96.5,58.5</position>
<gparam>LABEL_TEXT Seletores (S)</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>451</ID>
<type>AA_LABEL</type>
<position>31,73</position>
<gparam>LABEL_TEXT 74HC283</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>452</ID>
<type>AA_LABEL</type>
<position>22,73</position>
<gparam>LABEL_TEXT U4a</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>453</ID>
<type>AA_LABEL</type>
<position>40,73</position>
<gparam>LABEL_TEXT U4b</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>82</ID>
<type>AE_FULLADDER_4BIT</type>
<position>22,68</position>
<input>
<ID>IN_0</ID>46 </input>
<input>
<ID>IN_1</ID>45 </input>
<input>
<ID>IN_2</ID>44 </input>
<input>
<ID>IN_3</ID>43 </input>
<input>
<ID>IN_B_0</ID>102 </input>
<input>
<ID>IN_B_1</ID>103 </input>
<input>
<ID>IN_B_2</ID>104 </input>
<input>
<ID>IN_B_3</ID>105 </input>
<output>
<ID>OUT_0</ID>30 </output>
<output>
<ID>OUT_1</ID>31 </output>
<output>
<ID>OUT_2</ID>32 </output>
<output>
<ID>OUT_3</ID>33 </output>
<input>
<ID>carry_in</ID>42 </input>
<output>
<ID>carry_out</ID>51 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>84</ID>
<type>GA_LED</type>
<position>41.5,49</position>
<input>
<ID>N_in3</ID>26 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>86</ID>
<type>GA_LED</type>
<position>38.5,49</position>
<input>
<ID>N_in3</ID>27 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>88</ID>
<type>GA_LED</type>
<position>35.5,49</position>
<input>
<ID>N_in3</ID>28 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>90</ID>
<type>GA_LED</type>
<position>32.5,49</position>
<input>
<ID>N_in3</ID>29 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>92</ID>
<type>AE_FULLADDER_4BIT</type>
<position>40,68</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>49 </input>
<input>
<ID>IN_2</ID>48 </input>
<input>
<ID>IN_3</ID>47 </input>
<input>
<ID>IN_B_0</ID>82 </input>
<input>
<ID>IN_B_1</ID>85 </input>
<input>
<ID>IN_B_2</ID>100 </input>
<input>
<ID>IN_B_3</ID>101 </input>
<output>
<ID>OUT_0</ID>26 </output>
<output>
<ID>OUT_1</ID>27 </output>
<output>
<ID>OUT_2</ID>28 </output>
<output>
<ID>OUT_3</ID>29 </output>
<input>
<ID>carry_in</ID>64 </input>
<output>
<ID>carry_out</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>93</ID>
<type>AA_LABEL</type>
<position>20.5,46.5</position>
<gparam>LABEL_TEXT G7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>94</ID>
<type>AA_LABEL</type>
<position>23.5,46.5</position>
<gparam>LABEL_TEXT G6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>95</ID>
<type>AA_LABEL</type>
<position>26.5,46.5</position>
<gparam>LABEL_TEXT G5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>96</ID>
<type>AA_LABEL</type>
<position>29.5,46.5</position>
<gparam>LABEL_TEXT G4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>97</ID>
<type>GA_LED</type>
<position>29.5,49</position>
<input>
<ID>N_in3</ID>30 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>98</ID>
<type>GA_LED</type>
<position>26.5,49</position>
<input>
<ID>N_in3</ID>31 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>99</ID>
<type>GA_LED</type>
<position>23.5,49</position>
<input>
<ID>N_in3</ID>32 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>100</ID>
<type>GA_LED</type>
<position>20.5,49</position>
<input>
<ID>N_in3</ID>33 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>101</ID>
<type>AA_TOGGLE</type>
<position>17,143</position>
<output>
<ID>OUT_0</ID>43 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>102</ID>
<type>AA_TOGGLE</type>
<position>20,143</position>
<output>
<ID>OUT_0</ID>44 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>103</ID>
<type>AA_TOGGLE</type>
<position>23,143</position>
<output>
<ID>OUT_0</ID>45 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>104</ID>
<type>AA_TOGGLE</type>
<position>26,143</position>
<output>
<ID>OUT_0</ID>46 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>105</ID>
<type>AA_TOGGLE</type>
<position>29,143</position>
<output>
<ID>OUT_0</ID>47 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>106</ID>
<type>AA_TOGGLE</type>
<position>32,143</position>
<output>
<ID>OUT_0</ID>48 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>107</ID>
<type>AA_TOGGLE</type>
<position>35,143</position>
<output>
<ID>OUT_0</ID>49 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>108</ID>
<type>AA_TOGGLE</type>
<position>38,143</position>
<output>
<ID>OUT_0</ID>50 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>138</ID>
<type>AA_LABEL</type>
<position>16,46.5</position>
<gparam>LABEL_TEXT G8</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>139</ID>
<type>GA_LED</type>
<position>16,49</position>
<input>
<ID>N_in3</ID>51 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>148</ID>
<type>AA_TOGGLE</type>
<position>95,64</position>
<output>
<ID>OUT_0</ID>107 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>149</ID>
<type>AA_TOGGLE</type>
<position>98,64</position>
<output>
<ID>OUT_0</ID>106 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>150</ID>
<type>AA_TOGGLE</type>
<position>101,64</position>
<output>
<ID>OUT_0</ID>64 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>151</ID>
<type>AA_LABEL</type>
<position>95,61.5</position>
<gparam>LABEL_TEXT S2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>152</ID>
<type>AA_LABEL</type>
<position>98,61.5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>153</ID>
<type>AA_LABEL</type>
<position>101,61.5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>155</ID>
<type>AA_AND2</type>
<position>61,105</position>
<input>
<ID>IN_0</ID>106 </input>
<input>
<ID>IN_1</ID>91 </input>
<output>
<ID>OUT</ID>72 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>156</ID>
<type>AA_AND2</type>
<position>61,101</position>
<input>
<ID>IN_0</ID>107 </input>
<input>
<ID>IN_1</ID>90 </input>
<output>
<ID>OUT</ID>71 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>157</ID>
<type>AA_AND2</type>
<position>61,97</position>
<input>
<ID>IN_0</ID>106 </input>
<input>
<ID>IN_1</ID>89 </input>
<output>
<ID>OUT</ID>70 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>158</ID>
<type>AA_AND2</type>
<position>61,93</position>
<input>
<ID>IN_0</ID>107 </input>
<input>
<ID>IN_1</ID>88 </input>
<output>
<ID>OUT</ID>69 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>159</ID>
<type>AA_AND2</type>
<position>61,89</position>
<input>
<ID>IN_0</ID>106 </input>
<input>
<ID>IN_1</ID>87 </input>
<output>
<ID>OUT</ID>68 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>160</ID>
<type>AA_AND2</type>
<position>61,85</position>
<input>
<ID>IN_0</ID>107 </input>
<input>
<ID>IN_1</ID>86 </input>
<output>
<ID>OUT</ID>67 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>161</ID>
<type>AA_AND2</type>
<position>61,81</position>
<input>
<ID>IN_0</ID>106 </input>
<input>
<ID>IN_1</ID>83 </input>
<output>
<ID>OUT</ID>65 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>162</ID>
<type>AA_AND2</type>
<position>61,77</position>
<input>
<ID>IN_0</ID>107 </input>
<input>
<ID>IN_1</ID>84 </input>
<output>
<ID>OUT</ID>66 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>171</ID>
<type>AA_AND2</type>
<position>61,137</position>
<input>
<ID>IN_0</ID>106 </input>
<input>
<ID>IN_1</ID>95 </input>
<output>
<ID>OUT</ID>80 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>172</ID>
<type>AA_AND2</type>
<position>61,133</position>
<input>
<ID>IN_0</ID>107 </input>
<input>
<ID>IN_1</ID>99 </input>
<output>
<ID>OUT</ID>79 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>173</ID>
<type>AA_AND2</type>
<position>61,129</position>
<input>
<ID>IN_0</ID>106 </input>
<input>
<ID>IN_1</ID>94 </input>
<output>
<ID>OUT</ID>78 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>174</ID>
<type>AA_AND2</type>
<position>61,125</position>
<input>
<ID>IN_0</ID>107 </input>
<input>
<ID>IN_1</ID>98 </input>
<output>
<ID>OUT</ID>77 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>175</ID>
<type>AA_AND2</type>
<position>61,121</position>
<input>
<ID>IN_0</ID>106 </input>
<input>
<ID>IN_1</ID>93 </input>
<output>
<ID>OUT</ID>76 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>176</ID>
<type>AA_AND2</type>
<position>61,117</position>
<input>
<ID>IN_0</ID>107 </input>
<input>
<ID>IN_1</ID>96 </input>
<output>
<ID>OUT</ID>75 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>177</ID>
<type>AA_AND2</type>
<position>61,113</position>
<input>
<ID>IN_0</ID>106 </input>
<input>
<ID>IN_1</ID>92 </input>
<output>
<ID>OUT</ID>74 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>178</ID>
<type>AA_AND2</type>
<position>61,109</position>
<input>
<ID>IN_0</ID>107 </input>
<input>
<ID>IN_1</ID>97 </input>
<output>
<ID>OUT</ID>73 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>180</ID>
<type>AE_OR2</type>
<position>52.5,79</position>
<input>
<ID>IN_0</ID>66 </input>
<input>
<ID>IN_1</ID>65 </input>
<output>
<ID>OUT</ID>82 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>181</ID>
<type>AE_OR2</type>
<position>52.5,87</position>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>68 </input>
<output>
<ID>OUT</ID>85 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>182</ID>
<type>AE_OR2</type>
<position>52.5,95</position>
<input>
<ID>IN_0</ID>69 </input>
<input>
<ID>IN_1</ID>70 </input>
<output>
<ID>OUT</ID>100 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>183</ID>
<type>AE_OR2</type>
<position>52.5,103</position>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>72 </input>
<output>
<ID>OUT</ID>101 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>184</ID>
<type>AE_OR2</type>
<position>52.5,111</position>
<input>
<ID>IN_0</ID>73 </input>
<input>
<ID>IN_1</ID>74 </input>
<output>
<ID>OUT</ID>102 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>185</ID>
<type>AE_OR2</type>
<position>52.5,119</position>
<input>
<ID>IN_0</ID>75 </input>
<input>
<ID>IN_1</ID>76 </input>
<output>
<ID>OUT</ID>103 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>186</ID>
<type>AE_OR2</type>
<position>52.5,127</position>
<input>
<ID>IN_0</ID>77 </input>
<input>
<ID>IN_1</ID>78 </input>
<output>
<ID>OUT</ID>104 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>187</ID>
<type>AE_OR2</type>
<position>52.5,135</position>
<input>
<ID>IN_0</ID>79 </input>
<input>
<ID>IN_1</ID>80 </input>
<output>
<ID>OUT</ID>105 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>189</ID>
<type>AE_SMALL_INVERTER</type>
<position>69,78</position>
<input>
<ID>IN_0</ID>83 </input>
<output>
<ID>OUT_0</ID>84 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>190</ID>
<type>AE_SMALL_INVERTER</type>
<position>69,86</position>
<input>
<ID>IN_0</ID>87 </input>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>191</ID>
<type>AE_SMALL_INVERTER</type>
<position>69,94</position>
<input>
<ID>IN_0</ID>89 </input>
<output>
<ID>OUT_0</ID>88 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>192</ID>
<type>AE_SMALL_INVERTER</type>
<position>69,102</position>
<input>
<ID>IN_0</ID>91 </input>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41.5,50,41.5,64</points>
<connection>
<GID>92</GID>
<name>OUT_0</name></connection>
<connection>
<GID>84</GID>
<name>N_in3</name></connection></vsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,50,38.5,62</points>
<connection>
<GID>86</GID>
<name>N_in3</name></connection>
<intersection>62 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>40.5,62,40.5,64</points>
<connection>
<GID>92</GID>
<name>OUT_1</name></connection>
<intersection>62 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>38.5,62,40.5,62</points>
<intersection>38.5 0</intersection>
<intersection>40.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,50,35.5,63</points>
<connection>
<GID>88</GID>
<name>N_in3</name></connection>
<intersection>63 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>35.5,63,39.5,63</points>
<intersection>35.5 0</intersection>
<intersection>39.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>39.5,63,39.5,64</points>
<connection>
<GID>92</GID>
<name>OUT_2</name></connection>
<intersection>63 3</intersection></vsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,50,32.5,64</points>
<connection>
<GID>90</GID>
<name>N_in3</name></connection>
<intersection>64 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>32.5,64,38.5,64</points>
<connection>
<GID>92</GID>
<name>OUT_3</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,50,29.5,64</points>
<connection>
<GID>97</GID>
<name>N_in3</name></connection>
<intersection>64 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>23.5,64,29.5,64</points>
<connection>
<GID>82</GID>
<name>OUT_0</name></connection>
<intersection>29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,50,26.5,63</points>
<connection>
<GID>98</GID>
<name>N_in3</name></connection>
<intersection>63 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>22.5,63,26.5,63</points>
<intersection>22.5 4</intersection>
<intersection>26.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>22.5,63,22.5,64</points>
<connection>
<GID>82</GID>
<name>OUT_1</name></connection>
<intersection>63 3</intersection></vsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,62,21.5,64</points>
<connection>
<GID>82</GID>
<name>OUT_2</name></connection>
<intersection>62 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>21.5,62,23.5,62</points>
<intersection>21.5 0</intersection>
<intersection>23.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>23.5,50,23.5,62</points>
<connection>
<GID>99</GID>
<name>N_in3</name></connection>
<intersection>62 4</intersection></vsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,50,20.5,64</points>
<connection>
<GID>82</GID>
<name>OUT_3</name></connection>
<connection>
<GID>100</GID>
<name>N_in3</name></connection></vsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30,69,32,69</points>
<connection>
<GID>82</GID>
<name>carry_in</name></connection>
<connection>
<GID>92</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,72,17,141</points>
<connection>
<GID>82</GID>
<name>IN_3</name></connection>
<connection>
<GID>101</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,72,18,140</points>
<connection>
<GID>82</GID>
<name>IN_2</name></connection>
<intersection>140 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>20,140,20,141</points>
<connection>
<GID>102</GID>
<name>OUT_0</name></connection>
<intersection>140 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>18,140,20,140</points>
<intersection>18 0</intersection>
<intersection>20 1</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,72,19,139</points>
<connection>
<GID>82</GID>
<name>IN_1</name></connection>
<intersection>139 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>23,139,23,141</points>
<connection>
<GID>103</GID>
<name>OUT_0</name></connection>
<intersection>139 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>19,139,23,139</points>
<intersection>19 0</intersection>
<intersection>23 1</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,138,26,141</points>
<connection>
<GID>104</GID>
<name>OUT_0</name></connection>
<intersection>138 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>20,138,26,138</points>
<intersection>20 5</intersection>
<intersection>26 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>20,72,20,138</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<intersection>138 4</intersection></vsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,138,29,141</points>
<connection>
<GID>105</GID>
<name>OUT_0</name></connection>
<intersection>138 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>29,138,35,138</points>
<intersection>29 0</intersection>
<intersection>35 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>35,72,35,138</points>
<connection>
<GID>92</GID>
<name>IN_3</name></connection>
<intersection>138 3</intersection></vsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,72,36,139</points>
<connection>
<GID>92</GID>
<name>IN_2</name></connection>
<intersection>139 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>32,139,32,141</points>
<connection>
<GID>106</GID>
<name>OUT_0</name></connection>
<intersection>139 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>32,139,36,139</points>
<intersection>32 1</intersection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,72,37,140</points>
<connection>
<GID>92</GID>
<name>IN_1</name></connection>
<intersection>140 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>35,140,35,141</points>
<connection>
<GID>107</GID>
<name>OUT_0</name></connection>
<intersection>140 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>35,140,37,140</points>
<intersection>35 1</intersection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,72,38,141</points>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<connection>
<GID>108</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11.5,62,11.5,69</points>
<intersection>62 2</intersection>
<intersection>69 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>11.5,69,14,69</points>
<connection>
<GID>82</GID>
<name>carry_out</name></connection>
<intersection>11.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11.5,62,16,62</points>
<intersection>11.5 0</intersection>
<intersection>16 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>16,50,16,62</points>
<connection>
<GID>139</GID>
<name>N_in3</name></connection>
<intersection>62 2</intersection></vsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,66,101,69</points>
<connection>
<GID>150</GID>
<name>OUT_0</name></connection>
<intersection>69 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48,69,101,69</points>
<connection>
<GID>92</GID>
<name>carry_in</name></connection>
<intersection>101 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,80,56.5,81</points>
<intersection>80 2</intersection>
<intersection>81 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56.5,81,58,81</points>
<connection>
<GID>161</GID>
<name>OUT</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>55.5,80,56.5,80</points>
<connection>
<GID>180</GID>
<name>IN_1</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,77,56.5,78</points>
<intersection>77 2</intersection>
<intersection>78 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55.5,78,56.5,78</points>
<connection>
<GID>180</GID>
<name>IN_0</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,77,58,77</points>
<connection>
<GID>162</GID>
<name>OUT</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,85,56.5,86</points>
<intersection>85 2</intersection>
<intersection>86 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55.5,86,56.5,86</points>
<connection>
<GID>181</GID>
<name>IN_0</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,85,58,85</points>
<connection>
<GID>160</GID>
<name>OUT</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,88,56.5,89</points>
<intersection>88 1</intersection>
<intersection>89 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55.5,88,56.5,88</points>
<connection>
<GID>181</GID>
<name>IN_1</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,89,58,89</points>
<connection>
<GID>159</GID>
<name>OUT</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,93,56.5,94</points>
<intersection>93 2</intersection>
<intersection>94 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55.5,94,56.5,94</points>
<connection>
<GID>182</GID>
<name>IN_0</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,93,58,93</points>
<connection>
<GID>158</GID>
<name>OUT</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,96,56.5,97</points>
<intersection>96 1</intersection>
<intersection>97 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55.5,96,56.5,96</points>
<connection>
<GID>182</GID>
<name>IN_1</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,97,58,97</points>
<connection>
<GID>157</GID>
<name>OUT</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,101,56.5,102</points>
<intersection>101 2</intersection>
<intersection>102 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55.5,102,56.5,102</points>
<connection>
<GID>183</GID>
<name>IN_0</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,101,58,101</points>
<connection>
<GID>156</GID>
<name>OUT</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,104,56.5,105</points>
<intersection>104 1</intersection>
<intersection>105 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55.5,104,56.5,104</points>
<connection>
<GID>183</GID>
<name>IN_1</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,105,58,105</points>
<connection>
<GID>155</GID>
<name>OUT</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,109,56.5,110</points>
<intersection>109 2</intersection>
<intersection>110 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55.5,110,56.5,110</points>
<connection>
<GID>184</GID>
<name>IN_0</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,109,58,109</points>
<connection>
<GID>178</GID>
<name>OUT</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,112,56.5,113</points>
<intersection>112 1</intersection>
<intersection>113 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55.5,112,56.5,112</points>
<connection>
<GID>184</GID>
<name>IN_1</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,113,58,113</points>
<connection>
<GID>177</GID>
<name>OUT</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,117,56.5,118</points>
<intersection>117 2</intersection>
<intersection>118 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55.5,118,56.5,118</points>
<connection>
<GID>185</GID>
<name>IN_0</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,117,58,117</points>
<connection>
<GID>176</GID>
<name>OUT</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,120,56.5,121</points>
<intersection>120 1</intersection>
<intersection>121 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55.5,120,56.5,120</points>
<connection>
<GID>185</GID>
<name>IN_1</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,121,58,121</points>
<connection>
<GID>175</GID>
<name>OUT</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,125,56.5,126</points>
<intersection>125 2</intersection>
<intersection>126 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55.5,126,56.5,126</points>
<connection>
<GID>186</GID>
<name>IN_0</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,125,58,125</points>
<connection>
<GID>174</GID>
<name>OUT</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,128,56.5,129</points>
<intersection>128 1</intersection>
<intersection>129 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55.5,128,56.5,128</points>
<connection>
<GID>186</GID>
<name>IN_1</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,129,58,129</points>
<connection>
<GID>173</GID>
<name>OUT</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,133,56.5,134</points>
<intersection>133 2</intersection>
<intersection>134 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55.5,134,56.5,134</points>
<connection>
<GID>187</GID>
<name>IN_0</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,133,58,133</points>
<connection>
<GID>172</GID>
<name>OUT</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,136,56.5,137</points>
<intersection>136 1</intersection>
<intersection>137 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55.5,136,56.5,136</points>
<connection>
<GID>187</GID>
<name>IN_1</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,137,58,137</points>
<connection>
<GID>171</GID>
<name>OUT</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,72,45,79</points>
<connection>
<GID>92</GID>
<name>IN_B_0</name></connection>
<intersection>79 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,79,49.5,79</points>
<connection>
<GID>180</GID>
<name>OUT</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92,82,92,141</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<intersection>82 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64,82,92,82</points>
<connection>
<GID>161</GID>
<name>IN_1</name></connection>
<intersection>71 2</intersection>
<intersection>92 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71,78,71,82</points>
<connection>
<GID>189</GID>
<name>IN_0</name></connection>
<intersection>82 1</intersection></vsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64,78,67,78</points>
<connection>
<GID>162</GID>
<name>IN_1</name></connection>
<connection>
<GID>189</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,72,44,87</points>
<connection>
<GID>92</GID>
<name>IN_B_1</name></connection>
<intersection>87 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44,87,49.5,87</points>
<connection>
<GID>181</GID>
<name>OUT</name></connection>
<intersection>44 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64,86,67,86</points>
<connection>
<GID>160</GID>
<name>IN_1</name></connection>
<connection>
<GID>190</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,90,89,141</points>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection>
<intersection>90 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64,90,89,90</points>
<connection>
<GID>159</GID>
<name>IN_1</name></connection>
<intersection>71 2</intersection>
<intersection>89 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71,86,71,90</points>
<connection>
<GID>190</GID>
<name>IN_0</name></connection>
<intersection>90 1</intersection></vsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64,94,67,94</points>
<connection>
<GID>158</GID>
<name>IN_1</name></connection>
<connection>
<GID>191</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86,98,86,141</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<intersection>98 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64,98,86,98</points>
<connection>
<GID>157</GID>
<name>IN_1</name></connection>
<intersection>71 2</intersection>
<intersection>86 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71,94,71,98</points>
<connection>
<GID>191</GID>
<name>IN_0</name></connection>
<intersection>98 1</intersection></vsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64,102,67,102</points>
<connection>
<GID>156</GID>
<name>IN_1</name></connection>
<connection>
<GID>192</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83,106,83,141</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>106 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64,106,83,106</points>
<connection>
<GID>155</GID>
<name>IN_1</name></connection>
<intersection>71 2</intersection>
<intersection>83 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71,102,71,106</points>
<connection>
<GID>192</GID>
<name>IN_0</name></connection>
<intersection>106 1</intersection></vsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,114,80,141</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>114 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64,114,80,114</points>
<connection>
<GID>177</GID>
<name>IN_1</name></connection>
<intersection>71 2</intersection>
<intersection>80 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71,110,71,114</points>
<connection>
<GID>193</GID>
<name>IN_0</name></connection>
<intersection>114 1</intersection></vsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77,122,77,141</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<intersection>122 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64,122,77,122</points>
<connection>
<GID>175</GID>
<name>IN_1</name></connection>
<intersection>71 2</intersection>
<intersection>77 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71,118,71,122</points>
<connection>
<GID>194</GID>
<name>IN_0</name></connection>
<intersection>122 1</intersection></vsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74,130,74,141</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>130 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64,130,74,130</points>
<connection>
<GID>173</GID>
<name>IN_1</name></connection>
<intersection>71 2</intersection>
<intersection>74 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>71,126,71,130</points>
<connection>
<GID>195</GID>
<name>IN_0</name></connection>
<intersection>130 1</intersection></vsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71,134,71,141</points>
<connection>
<GID>196</GID>
<name>IN_0</name></connection>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection>
<intersection>138 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64,138,71,138</points>
<connection>
<GID>171</GID>
<name>IN_1</name></connection>
<intersection>71 0</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64,118,67,118</points>
<connection>
<GID>176</GID>
<name>IN_1</name></connection>
<connection>
<GID>194</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64,110,67,110</points>
<connection>
<GID>178</GID>
<name>IN_1</name></connection>
<connection>
<GID>193</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64,126,67,126</points>
<connection>
<GID>174</GID>
<name>IN_1</name></connection>
<connection>
<GID>195</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64,134,67,134</points>
<connection>
<GID>172</GID>
<name>IN_1</name></connection>
<connection>
<GID>196</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43,72,43,95</points>
<connection>
<GID>92</GID>
<name>IN_B_2</name></connection>
<intersection>95 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43,95,49.5,95</points>
<connection>
<GID>182</GID>
<name>OUT</name></connection>
<intersection>43 0</intersection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42,72,42,103</points>
<connection>
<GID>92</GID>
<name>IN_B_3</name></connection>
<intersection>103 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42,103,49.5,103</points>
<connection>
<GID>183</GID>
<name>OUT</name></connection>
<intersection>42 0</intersection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,72,27,111</points>
<connection>
<GID>82</GID>
<name>IN_B_0</name></connection>
<intersection>111 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,111,49.5,111</points>
<connection>
<GID>184</GID>
<name>OUT</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,72,26,119</points>
<connection>
<GID>82</GID>
<name>IN_B_1</name></connection>
<intersection>119 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,119,49.5,119</points>
<connection>
<GID>185</GID>
<name>OUT</name></connection>
<intersection>26 0</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,72,25,127</points>
<connection>
<GID>82</GID>
<name>IN_B_2</name></connection>
<intersection>127 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,127,49.5,127</points>
<connection>
<GID>186</GID>
<name>OUT</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,72,24,135</points>
<connection>
<GID>82</GID>
<name>IN_B_3</name></connection>
<intersection>135 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24,135,49.5,135</points>
<connection>
<GID>187</GID>
<name>OUT</name></connection>
<intersection>24 0</intersection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98,66,98,136</points>
<connection>
<GID>149</GID>
<name>OUT_0</name></connection>
<intersection>80 1</intersection>
<intersection>88 3</intersection>
<intersection>96 5</intersection>
<intersection>104 7</intersection>
<intersection>112 9</intersection>
<intersection>120 11</intersection>
<intersection>128 13</intersection>
<intersection>136 15</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64,80,98,80</points>
<connection>
<GID>161</GID>
<name>IN_0</name></connection>
<intersection>98 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>64,88,98,88</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<intersection>98 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>64,96,98,96</points>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<intersection>98 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>64,104,98,104</points>
<connection>
<GID>155</GID>
<name>IN_0</name></connection>
<intersection>98 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>64,112,98,112</points>
<connection>
<GID>177</GID>
<name>IN_0</name></connection>
<intersection>98 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>64,120,98,120</points>
<connection>
<GID>175</GID>
<name>IN_0</name></connection>
<intersection>98 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>64,128,98,128</points>
<connection>
<GID>173</GID>
<name>IN_0</name></connection>
<intersection>98 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>64,136,98,136</points>
<connection>
<GID>171</GID>
<name>IN_0</name></connection>
<intersection>98 0</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95,66,95,132</points>
<connection>
<GID>148</GID>
<name>OUT_0</name></connection>
<intersection>76 1</intersection>
<intersection>84 3</intersection>
<intersection>92 5</intersection>
<intersection>100 7</intersection>
<intersection>108 9</intersection>
<intersection>116 11</intersection>
<intersection>124 13</intersection>
<intersection>132 15</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64,76,95,76</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>64,84,95,84</points>
<connection>
<GID>160</GID>
<name>IN_0</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>64,92,95,92</points>
<connection>
<GID>158</GID>
<name>IN_0</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>64,100,95,100</points>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>64,108,95,108</points>
<connection>
<GID>178</GID>
<name>IN_0</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>64,116,95,116</points>
<connection>
<GID>176</GID>
<name>IN_0</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>64,124,95,124</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>64,132,95,132</points>
<connection>
<GID>172</GID>
<name>IN_0</name></connection>
<intersection>95 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-67.1379,13.0412,226.438,-138.37</PageViewport>
<gate>
<ID>203</ID>
<type>AA_TOGGLE</type>
<position>109,-5</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>204</ID>
<type>AA_LABEL</type>
<position>109,-2.5</position>
<gparam>LABEL_TEXT S3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>205</ID>
<type>AA_TOGGLE</type>
<position>40,-5</position>
<output>
<ID>OUT_0</ID>235 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>206</ID>
<type>AA_TOGGLE</type>
<position>43,-5</position>
<output>
<ID>OUT_0</ID>237 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>207</ID>
<type>AA_TOGGLE</type>
<position>46,-5</position>
<output>
<ID>OUT_0</ID>239 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>208</ID>
<type>AA_TOGGLE</type>
<position>49,-5</position>
<output>
<ID>OUT_0</ID>241 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>209</ID>
<type>AA_TOGGLE</type>
<position>52,-5</position>
<output>
<ID>OUT_0</ID>243 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>210</ID>
<type>AA_TOGGLE</type>
<position>55,-5</position>
<output>
<ID>OUT_0</ID>245 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>211</ID>
<type>AA_TOGGLE</type>
<position>58,-5</position>
<output>
<ID>OUT_0</ID>247 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>212</ID>
<type>AA_TOGGLE</type>
<position>61,-5</position>
<output>
<ID>OUT_0</ID>249 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>213</ID>
<type>AA_LABEL</type>
<position>10,-2.5</position>
<gparam>LABEL_TEXT X7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>214</ID>
<type>AA_LABEL</type>
<position>13,-2.5</position>
<gparam>LABEL_TEXT X6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>407</ID>
<type>AA_LABEL</type>
<position>64.5,11.5</position>
<gparam>LABEL_TEXT Unidade Logica</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>215</ID>
<type>AA_LABEL</type>
<position>16,-2.5</position>
<gparam>LABEL_TEXT X5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>216</ID>
<type>AA_LABEL</type>
<position>19,-2.5</position>
<gparam>LABEL_TEXT X4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>217</ID>
<type>AA_LABEL</type>
<position>22,-2.5</position>
<gparam>LABEL_TEXT X3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>218</ID>
<type>AA_LABEL</type>
<position>25,-2.5</position>
<gparam>LABEL_TEXT X2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>219</ID>
<type>AA_LABEL</type>
<position>28,-2.5</position>
<gparam>LABEL_TEXT X1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>220</ID>
<type>AA_LABEL</type>
<position>31,-2.5</position>
<gparam>LABEL_TEXT X0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>221</ID>
<type>AA_LABEL</type>
<position>40,-2.5</position>
<gparam>LABEL_TEXT Y7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>222</ID>
<type>AA_LABEL</type>
<position>43,-2.5</position>
<gparam>LABEL_TEXT Y6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>223</ID>
<type>AA_LABEL</type>
<position>46,-2.5</position>
<gparam>LABEL_TEXT Y5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>224</ID>
<type>AA_LABEL</type>
<position>49,-2.5</position>
<gparam>LABEL_TEXT Y4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>225</ID>
<type>AA_LABEL</type>
<position>52,-2.5</position>
<gparam>LABEL_TEXT Y3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>226</ID>
<type>AA_LABEL</type>
<position>55,-2.5</position>
<gparam>LABEL_TEXT Y2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>227</ID>
<type>AA_LABEL</type>
<position>58,-2.5</position>
<gparam>LABEL_TEXT Y1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>228</ID>
<type>AA_LABEL</type>
<position>61,-2.5</position>
<gparam>LABEL_TEXT Y0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>229</ID>
<type>AA_LABEL</type>
<position>132.5,-75</position>
<gparam>LABEL_TEXT G3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>230</ID>
<type>AA_LABEL</type>
<position>132.5,-79</position>
<gparam>LABEL_TEXT G2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>231</ID>
<type>AA_LABEL</type>
<position>132.5,-83</position>
<gparam>LABEL_TEXT G1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>232</ID>
<type>AA_LABEL</type>
<position>132.5,-86.5</position>
<gparam>LABEL_TEXT G0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>234</ID>
<type>GA_LED</type>
<position>130,-59</position>
<input>
<ID>N_in0</ID>224 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>235</ID>
<type>GA_LED</type>
<position>130,-63</position>
<input>
<ID>N_in0</ID>225 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>236</ID>
<type>GA_LED</type>
<position>130,-67</position>
<input>
<ID>N_in0</ID>226 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>237</ID>
<type>GA_LED</type>
<position>130,-71</position>
<input>
<ID>N_in0</ID>227 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>239</ID>
<type>AA_LABEL</type>
<position>132.5,-59</position>
<gparam>LABEL_TEXT G7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>240</ID>
<type>AA_LABEL</type>
<position>132.5,-63</position>
<gparam>LABEL_TEXT G6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>241</ID>
<type>AA_LABEL</type>
<position>132.5,-67</position>
<gparam>LABEL_TEXT G5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>242</ID>
<type>AA_LABEL</type>
<position>132.5,-71</position>
<gparam>LABEL_TEXT G4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>243</ID>
<type>GA_LED</type>
<position>130,-75</position>
<input>
<ID>N_in0</ID>228 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>244</ID>
<type>GA_LED</type>
<position>130,-79</position>
<input>
<ID>N_in0</ID>229 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>245</ID>
<type>GA_LED</type>
<position>130,-83</position>
<input>
<ID>N_in0</ID>230 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>246</ID>
<type>GA_LED</type>
<position>130,-87</position>
<input>
<ID>N_in0</ID>231 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>247</ID>
<type>AA_TOGGLE</type>
<position>10,-5</position>
<output>
<ID>OUT_0</ID>236 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>248</ID>
<type>AA_TOGGLE</type>
<position>13,-5</position>
<output>
<ID>OUT_0</ID>238 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>249</ID>
<type>AA_TOGGLE</type>
<position>16,-5</position>
<output>
<ID>OUT_0</ID>240 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>250</ID>
<type>AA_TOGGLE</type>
<position>19,-5</position>
<output>
<ID>OUT_0</ID>242 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>251</ID>
<type>AA_TOGGLE</type>
<position>21.5,-5</position>
<output>
<ID>OUT_0</ID>244 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>252</ID>
<type>AA_TOGGLE</type>
<position>25,-5</position>
<output>
<ID>OUT_0</ID>246 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>253</ID>
<type>AA_TOGGLE</type>
<position>28,-5</position>
<output>
<ID>OUT_0</ID>248 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>254</ID>
<type>AA_TOGGLE</type>
<position>31,-5</position>
<output>
<ID>OUT_0</ID>250 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>257</ID>
<type>AA_TOGGLE</type>
<position>112,-5</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>258</ID>
<type>AA_TOGGLE</type>
<position>115,-5</position>
<output>
<ID>OUT_0</ID>223 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>259</ID>
<type>AA_TOGGLE</type>
<position>118,-5</position>
<output>
<ID>OUT_0</ID>222 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>260</ID>
<type>AA_LABEL</type>
<position>112,-2.5</position>
<gparam>LABEL_TEXT S2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>261</ID>
<type>AA_LABEL</type>
<position>115,-2.5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>454</ID>
<type>AA_LABEL</type>
<position>20.5,1</position>
<gparam>LABEL_TEXT Entradas (X)</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>262</ID>
<type>AA_LABEL</type>
<position>118,-2.5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>455</ID>
<type>AA_LABEL</type>
<position>50.5,1</position>
<gparam>LABEL_TEXT Entradas (Y)</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>456</ID>
<type>AA_LABEL</type>
<position>113.5,1</position>
<gparam>LABEL_TEXT Seletores (S)</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>457</ID>
<type>AA_LABEL</type>
<position>142.5,-72.5</position>
<gparam>LABEL_TEXT Saidas (G)</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>458</ID>
<type>AA_LABEL</type>
<position>67,-11</position>
<gparam>LABEL_TEXT 74HC08</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>460</ID>
<type>AA_LABEL</type>
<position>67,-45</position>
<gparam>LABEL_TEXT 74HC32</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>461</ID>
<type>AA_LABEL</type>
<position>67,-79</position>
<gparam>LABEL_TEXT 74HC86</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>462</ID>
<type>AA_LABEL</type>
<position>67,-114</position>
<gparam>LABEL_TEXT 74HC04</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>463</ID>
<type>AA_LABEL</type>
<position>62.5,-14</position>
<gparam>LABEL_TEXT U1a</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>464</ID>
<type>AA_LABEL</type>
<position>62.5,-18</position>
<gparam>LABEL_TEXT U1b</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>465</ID>
<type>AA_LABEL</type>
<position>62.5,-22</position>
<gparam>LABEL_TEXT U1c</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>466</ID>
<type>AA_LABEL</type>
<position>62.5,-26</position>
<gparam>LABEL_TEXT U1d</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>467</ID>
<type>AA_LABEL</type>
<position>62.5,-30</position>
<gparam>LABEL_TEXT U1e</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>468</ID>
<type>AA_LABEL</type>
<position>62.5,-34</position>
<gparam>LABEL_TEXT U1f</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>469</ID>
<type>AA_LABEL</type>
<position>62.5,-38</position>
<gparam>LABEL_TEXT U1g</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>470</ID>
<type>AA_LABEL</type>
<position>62.5,-42</position>
<gparam>LABEL_TEXT U1h</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>471</ID>
<type>AA_LABEL</type>
<position>62.5,-48</position>
<gparam>LABEL_TEXT U2a</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>472</ID>
<type>AA_LABEL</type>
<position>62.5,-52</position>
<gparam>LABEL_TEXT U2b</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>473</ID>
<type>AA_LABEL</type>
<position>62.5,-56</position>
<gparam>LABEL_TEXT U2c</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>474</ID>
<type>AA_LABEL</type>
<position>62.5,-60</position>
<gparam>LABEL_TEXT U2d</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>475</ID>
<type>AA_LABEL</type>
<position>62.5,-64</position>
<gparam>LABEL_TEXT U2e</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>476</ID>
<type>AA_LABEL</type>
<position>62.5,-68</position>
<gparam>LABEL_TEXT U2f</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>477</ID>
<type>AA_LABEL</type>
<position>62.5,-72</position>
<gparam>LABEL_TEXT U2g</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>478</ID>
<type>AA_LABEL</type>
<position>62.5,-76</position>
<gparam>LABEL_TEXT U2h</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>479</ID>
<type>AA_LABEL</type>
<position>62.5,-82</position>
<gparam>LABEL_TEXT U3a</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>480</ID>
<type>AA_LABEL</type>
<position>62.5,-86</position>
<gparam>LABEL_TEXT U3b</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>481</ID>
<type>AA_LABEL</type>
<position>62.5,-90</position>
<gparam>LABEL_TEXT U3c</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>482</ID>
<type>AA_LABEL</type>
<position>62.5,-94</position>
<gparam>LABEL_TEXT U3d</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>483</ID>
<type>AA_LABEL</type>
<position>62.5,-98</position>
<gparam>LABEL_TEXT U3e</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>484</ID>
<type>AA_LABEL</type>
<position>62.5,-102</position>
<gparam>LABEL_TEXT U3f</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>292</ID>
<type>AA_AND2</type>
<position>67,-14</position>
<input>
<ID>IN_0</ID>235 </input>
<input>
<ID>IN_1</ID>236 </input>
<output>
<ID>OUT</ID>213 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>485</ID>
<type>AA_LABEL</type>
<position>62.5,-106</position>
<gparam>LABEL_TEXT U3g</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>293</ID>
<type>AA_AND2</type>
<position>67,-18</position>
<input>
<ID>IN_0</ID>237 </input>
<input>
<ID>IN_1</ID>238 </input>
<output>
<ID>OUT</ID>221 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>486</ID>
<type>AA_LABEL</type>
<position>62.5,-110</position>
<gparam>LABEL_TEXT U3h</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>294</ID>
<type>AA_AND2</type>
<position>67,-22</position>
<input>
<ID>IN_0</ID>239 </input>
<input>
<ID>IN_1</ID>240 </input>
<output>
<ID>OUT</ID>220 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>487</ID>
<type>AA_LABEL</type>
<position>63,-116.5</position>
<gparam>LABEL_TEXT U4a</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>295</ID>
<type>AA_AND2</type>
<position>67,-26</position>
<input>
<ID>IN_0</ID>241 </input>
<input>
<ID>IN_1</ID>242 </input>
<output>
<ID>OUT</ID>218 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>488</ID>
<type>AA_LABEL</type>
<position>63,-119.5</position>
<gparam>LABEL_TEXT U4b</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>296</ID>
<type>AA_AND2</type>
<position>67,-30</position>
<input>
<ID>IN_0</ID>243 </input>
<input>
<ID>IN_1</ID>244 </input>
<output>
<ID>OUT</ID>217 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>489</ID>
<type>AA_LABEL</type>
<position>63,-122.5</position>
<gparam>LABEL_TEXT U4c</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>297</ID>
<type>AA_AND2</type>
<position>67,-34</position>
<input>
<ID>IN_0</ID>245 </input>
<input>
<ID>IN_1</ID>246 </input>
<output>
<ID>OUT</ID>216 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>490</ID>
<type>AA_LABEL</type>
<position>63,-125.5</position>
<gparam>LABEL_TEXT U4d</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>298</ID>
<type>AA_AND2</type>
<position>67,-38</position>
<input>
<ID>IN_0</ID>247 </input>
<input>
<ID>IN_1</ID>248 </input>
<output>
<ID>OUT</ID>215 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>491</ID>
<type>AA_LABEL</type>
<position>63,-128.5</position>
<gparam>LABEL_TEXT U4e</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>299</ID>
<type>AA_AND2</type>
<position>67,-42</position>
<input>
<ID>IN_0</ID>249 </input>
<input>
<ID>IN_1</ID>250 </input>
<output>
<ID>OUT</ID>214 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>492</ID>
<type>AA_LABEL</type>
<position>63,-131.5</position>
<gparam>LABEL_TEXT U4f</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>493</ID>
<type>AA_LABEL</type>
<position>63,-134.5</position>
<gparam>LABEL_TEXT U4g</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>301</ID>
<type>AE_OR2</type>
<position>67,-48</position>
<input>
<ID>IN_0</ID>235 </input>
<input>
<ID>IN_1</ID>236 </input>
<output>
<ID>OUT</ID>212 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>494</ID>
<type>AA_LABEL</type>
<position>63,-137.5</position>
<gparam>LABEL_TEXT U4h</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>302</ID>
<type>AE_OR2</type>
<position>67,-52</position>
<input>
<ID>IN_0</ID>237 </input>
<input>
<ID>IN_1</ID>238 </input>
<output>
<ID>OUT</ID>211 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>303</ID>
<type>AE_OR2</type>
<position>67,-56</position>
<input>
<ID>IN_0</ID>239 </input>
<input>
<ID>IN_1</ID>240 </input>
<output>
<ID>OUT</ID>210 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>304</ID>
<type>AE_OR2</type>
<position>67,-60</position>
<input>
<ID>IN_0</ID>241 </input>
<input>
<ID>IN_1</ID>242 </input>
<output>
<ID>OUT</ID>209 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>305</ID>
<type>AE_OR2</type>
<position>67,-64</position>
<input>
<ID>IN_0</ID>243 </input>
<input>
<ID>IN_1</ID>244 </input>
<output>
<ID>OUT</ID>208 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>306</ID>
<type>AE_OR2</type>
<position>67,-68</position>
<input>
<ID>IN_0</ID>245 </input>
<input>
<ID>IN_1</ID>246 </input>
<output>
<ID>OUT</ID>207 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>307</ID>
<type>AE_OR2</type>
<position>67,-72</position>
<input>
<ID>IN_0</ID>247 </input>
<input>
<ID>IN_1</ID>248 </input>
<output>
<ID>OUT</ID>206 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>308</ID>
<type>AE_OR2</type>
<position>67,-76</position>
<input>
<ID>IN_0</ID>249 </input>
<input>
<ID>IN_1</ID>250 </input>
<output>
<ID>OUT</ID>205 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>310</ID>
<type>AI_XOR2</type>
<position>67.5,-82</position>
<input>
<ID>IN_0</ID>235 </input>
<input>
<ID>IN_1</ID>236 </input>
<output>
<ID>OUT</ID>197 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>503</ID>
<type>AA_LABEL</type>
<position>107,-16</position>
<gparam>LABEL_TEXT 74LS253</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>311</ID>
<type>AI_XOR2</type>
<position>67.5,-86</position>
<input>
<ID>IN_0</ID>237 </input>
<input>
<ID>IN_1</ID>238 </input>
<output>
<ID>OUT</ID>204 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>504</ID>
<type>AA_LABEL</type>
<position>107,-29</position>
<gparam>LABEL_TEXT U5a</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>312</ID>
<type>AI_XOR2</type>
<position>67.5,-90</position>
<input>
<ID>IN_0</ID>239 </input>
<input>
<ID>IN_1</ID>240 </input>
<output>
<ID>OUT</ID>203 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>505</ID>
<type>AA_LABEL</type>
<position>107,-43</position>
<gparam>LABEL_TEXT U5b</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>313</ID>
<type>AI_XOR2</type>
<position>67.5,-94</position>
<input>
<ID>IN_0</ID>241 </input>
<input>
<ID>IN_1</ID>242 </input>
<output>
<ID>OUT</ID>202 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>506</ID>
<type>AA_LABEL</type>
<position>107,-57</position>
<gparam>LABEL_TEXT U5c</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>314</ID>
<type>AI_XOR2</type>
<position>67.5,-98</position>
<input>
<ID>IN_0</ID>243 </input>
<input>
<ID>IN_1</ID>244 </input>
<output>
<ID>OUT</ID>201 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>507</ID>
<type>AA_LABEL</type>
<position>107,-71</position>
<gparam>LABEL_TEXT U5d</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>315</ID>
<type>AI_XOR2</type>
<position>67.5,-102</position>
<input>
<ID>IN_0</ID>245 </input>
<input>
<ID>IN_1</ID>246 </input>
<output>
<ID>OUT</ID>200 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>508</ID>
<type>AA_LABEL</type>
<position>107,-85</position>
<gparam>LABEL_TEXT U5e</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>316</ID>
<type>AI_XOR2</type>
<position>67.5,-106</position>
<input>
<ID>IN_0</ID>247 </input>
<input>
<ID>IN_1</ID>248 </input>
<output>
<ID>OUT</ID>199 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>509</ID>
<type>AA_LABEL</type>
<position>107,-99</position>
<gparam>LABEL_TEXT U5f</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>317</ID>
<type>AI_XOR2</type>
<position>67.5,-110</position>
<input>
<ID>IN_0</ID>249 </input>
<input>
<ID>IN_1</ID>250 </input>
<output>
<ID>OUT</ID>198 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>510</ID>
<type>AA_LABEL</type>
<position>107,-113</position>
<gparam>LABEL_TEXT U5g</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>511</ID>
<type>AA_LABEL</type>
<position>107,-127</position>
<gparam>LABEL_TEXT U5h</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>323</ID>
<type>AE_SMALL_INVERTER</type>
<position>67,-116</position>
<input>
<ID>IN_0</ID>236 </input>
<output>
<ID>OUT_0</ID>189 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>324</ID>
<type>AE_SMALL_INVERTER</type>
<position>67,-119</position>
<input>
<ID>IN_0</ID>238 </input>
<output>
<ID>OUT_0</ID>190 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>325</ID>
<type>AE_SMALL_INVERTER</type>
<position>67,-122</position>
<input>
<ID>IN_0</ID>240 </input>
<output>
<ID>OUT_0</ID>191 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>326</ID>
<type>AE_SMALL_INVERTER</type>
<position>67,-125</position>
<input>
<ID>IN_0</ID>242 </input>
<output>
<ID>OUT_0</ID>192 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>327</ID>
<type>AE_SMALL_INVERTER</type>
<position>67,-128</position>
<input>
<ID>IN_0</ID>244 </input>
<output>
<ID>OUT_0</ID>193 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>328</ID>
<type>AE_SMALL_INVERTER</type>
<position>67,-131</position>
<input>
<ID>IN_0</ID>246 </input>
<output>
<ID>OUT_0</ID>194 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>329</ID>
<type>AE_SMALL_INVERTER</type>
<position>67,-134</position>
<input>
<ID>IN_0</ID>248 </input>
<output>
<ID>OUT_0</ID>195 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>330</ID>
<type>AE_SMALL_INVERTER</type>
<position>67,-137</position>
<input>
<ID>IN_0</ID>250 </input>
<output>
<ID>OUT_0</ID>196 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>332</ID>
<type>AE_MUX_4x1</type>
<position>107,-24</position>
<input>
<ID>IN_0</ID>213 </input>
<input>
<ID>IN_1</ID>212 </input>
<input>
<ID>IN_2</ID>197 </input>
<input>
<ID>IN_3</ID>189 </input>
<output>
<ID>OUT</ID>224 </output>
<input>
<ID>SEL_0</ID>222 </input>
<input>
<ID>SEL_1</ID>223 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>333</ID>
<type>AE_MUX_4x1</type>
<position>107,-38</position>
<input>
<ID>IN_0</ID>221 </input>
<input>
<ID>IN_1</ID>211 </input>
<input>
<ID>IN_2</ID>204 </input>
<input>
<ID>IN_3</ID>190 </input>
<output>
<ID>OUT</ID>225 </output>
<input>
<ID>SEL_0</ID>222 </input>
<input>
<ID>SEL_1</ID>223 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>334</ID>
<type>AE_MUX_4x1</type>
<position>107,-52</position>
<input>
<ID>IN_0</ID>220 </input>
<input>
<ID>IN_1</ID>210 </input>
<input>
<ID>IN_2</ID>203 </input>
<input>
<ID>IN_3</ID>191 </input>
<output>
<ID>OUT</ID>226 </output>
<input>
<ID>SEL_0</ID>222 </input>
<input>
<ID>SEL_1</ID>223 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>335</ID>
<type>AE_MUX_4x1</type>
<position>107,-66</position>
<input>
<ID>IN_0</ID>218 </input>
<input>
<ID>IN_1</ID>209 </input>
<input>
<ID>IN_2</ID>202 </input>
<input>
<ID>IN_3</ID>192 </input>
<output>
<ID>OUT</ID>227 </output>
<input>
<ID>SEL_0</ID>222 </input>
<input>
<ID>SEL_1</ID>223 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>336</ID>
<type>AE_MUX_4x1</type>
<position>107,-80</position>
<input>
<ID>IN_0</ID>217 </input>
<input>
<ID>IN_1</ID>208 </input>
<input>
<ID>IN_2</ID>201 </input>
<input>
<ID>IN_3</ID>193 </input>
<output>
<ID>OUT</ID>228 </output>
<input>
<ID>SEL_0</ID>222 </input>
<input>
<ID>SEL_1</ID>223 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>337</ID>
<type>AE_MUX_4x1</type>
<position>107,-94</position>
<input>
<ID>IN_0</ID>216 </input>
<input>
<ID>IN_1</ID>207 </input>
<input>
<ID>IN_2</ID>200 </input>
<input>
<ID>IN_3</ID>194 </input>
<output>
<ID>OUT</ID>229 </output>
<input>
<ID>SEL_0</ID>222 </input>
<input>
<ID>SEL_1</ID>223 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>338</ID>
<type>AE_MUX_4x1</type>
<position>107,-108</position>
<input>
<ID>IN_0</ID>215 </input>
<input>
<ID>IN_1</ID>206 </input>
<input>
<ID>IN_2</ID>199 </input>
<input>
<ID>IN_3</ID>195 </input>
<output>
<ID>OUT</ID>230 </output>
<input>
<ID>SEL_0</ID>222 </input>
<input>
<ID>SEL_1</ID>223 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>339</ID>
<type>AE_MUX_4x1</type>
<position>107,-122</position>
<input>
<ID>IN_0</ID>214 </input>
<input>
<ID>IN_1</ID>205 </input>
<input>
<ID>IN_2</ID>198 </input>
<input>
<ID>IN_3</ID>196 </input>
<output>
<ID>OUT</ID>231 </output>
<input>
<ID>SEL_0</ID>222 </input>
<input>
<ID>SEL_1</ID>223 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<wire>
<ID>193</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97,-128,97,-77</points>
<intersection>-128 2</intersection>
<intersection>-77 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>97,-77,104,-77</points>
<connection>
<GID>336</GID>
<name>IN_3</name></connection>
<intersection>97 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69,-128,97,-128</points>
<connection>
<GID>327</GID>
<name>OUT_0</name></connection>
<intersection>97 0</intersection></hsegment></shape></wire>
<wire>
<ID>194</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98,-131,98,-91</points>
<intersection>-131 2</intersection>
<intersection>-91 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98,-91,104,-91</points>
<connection>
<GID>337</GID>
<name>IN_3</name></connection>
<intersection>98 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69,-131,98,-131</points>
<connection>
<GID>328</GID>
<name>OUT_0</name></connection>
<intersection>98 0</intersection></hsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-134,99,-105</points>
<intersection>-134 2</intersection>
<intersection>-105 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99,-105,104,-105</points>
<connection>
<GID>338</GID>
<name>IN_3</name></connection>
<intersection>99 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69,-134,99,-134</points>
<connection>
<GID>329</GID>
<name>OUT_0</name></connection>
<intersection>99 0</intersection></hsegment></shape></wire>
<wire>
<ID>196</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-137,100,-119</points>
<intersection>-137 2</intersection>
<intersection>-119 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100,-119,104,-119</points>
<connection>
<GID>339</GID>
<name>IN_3</name></connection>
<intersection>100 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69,-137,100,-137</points>
<connection>
<GID>330</GID>
<name>OUT_0</name></connection>
<intersection>100 0</intersection></hsegment></shape></wire>
<wire>
<ID>197</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,-82,85,-23</points>
<intersection>-82 2</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85,-23,104,-23</points>
<connection>
<GID>332</GID>
<name>IN_2</name></connection>
<intersection>85 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70.5,-82,85,-82</points>
<connection>
<GID>310</GID>
<name>OUT</name></connection>
<intersection>85 0</intersection></hsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-121,90,-110</points>
<intersection>-121 1</intersection>
<intersection>-110 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>90,-121,104,-121</points>
<connection>
<GID>339</GID>
<name>IN_2</name></connection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70.5,-110,90,-110</points>
<connection>
<GID>317</GID>
<name>OUT</name></connection>
<intersection>90 0</intersection></hsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-107,90,-106</points>
<intersection>-107 1</intersection>
<intersection>-106 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>90,-107,104,-107</points>
<connection>
<GID>338</GID>
<name>IN_2</name></connection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70.5,-106,90,-106</points>
<connection>
<GID>316</GID>
<name>OUT</name></connection>
<intersection>90 0</intersection></hsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-102,90,-93</points>
<intersection>-102 2</intersection>
<intersection>-93 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>90,-93,104,-93</points>
<connection>
<GID>337</GID>
<name>IN_2</name></connection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70.5,-102,90,-102</points>
<connection>
<GID>315</GID>
<name>OUT</name></connection>
<intersection>90 0</intersection></hsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,-98,89,-79</points>
<intersection>-98 2</intersection>
<intersection>-79 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>89,-79,104,-79</points>
<connection>
<GID>336</GID>
<name>IN_2</name></connection>
<intersection>89 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70.5,-98,89,-98</points>
<connection>
<GID>314</GID>
<name>OUT</name></connection>
<intersection>89 0</intersection></hsegment></shape></wire>
<wire>
<ID>202</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,-94,88,-65</points>
<intersection>-94 2</intersection>
<intersection>-65 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>88,-65,104,-65</points>
<connection>
<GID>335</GID>
<name>IN_2</name></connection>
<intersection>88 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70.5,-94,88,-94</points>
<connection>
<GID>313</GID>
<name>OUT</name></connection>
<intersection>88 0</intersection></hsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87,-90,87,-51</points>
<intersection>-90 2</intersection>
<intersection>-51 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>87,-51,104,-51</points>
<connection>
<GID>334</GID>
<name>IN_2</name></connection>
<intersection>87 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70.5,-90,87,-90</points>
<connection>
<GID>312</GID>
<name>OUT</name></connection>
<intersection>87 0</intersection></hsegment></shape></wire>
<wire>
<ID>204</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86,-86,86,-37</points>
<intersection>-86 2</intersection>
<intersection>-37 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>86,-37,104,-37</points>
<connection>
<GID>333</GID>
<name>IN_2</name></connection>
<intersection>86 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70.5,-86,86,-86</points>
<connection>
<GID>311</GID>
<name>OUT</name></connection>
<intersection>86 0</intersection></hsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78,-123,78,-76</points>
<intersection>-123 1</intersection>
<intersection>-76 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>78,-123,104,-123</points>
<connection>
<GID>339</GID>
<name>IN_1</name></connection>
<intersection>78 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70,-76,78,-76</points>
<connection>
<GID>308</GID>
<name>OUT</name></connection>
<intersection>78 0</intersection></hsegment></shape></wire>
<wire>
<ID>206</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79,-109,79,-72</points>
<intersection>-109 1</intersection>
<intersection>-72 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>79,-109,104,-109</points>
<connection>
<GID>338</GID>
<name>IN_1</name></connection>
<intersection>79 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70,-72,79,-72</points>
<connection>
<GID>307</GID>
<name>OUT</name></connection>
<intersection>79 0</intersection></hsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-95,80,-68</points>
<intersection>-95 1</intersection>
<intersection>-68 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80,-95,104,-95</points>
<connection>
<GID>337</GID>
<name>IN_1</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70,-68,80,-68</points>
<connection>
<GID>306</GID>
<name>OUT</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>208</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,-81,81,-64</points>
<intersection>-81 1</intersection>
<intersection>-64 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>81,-81,104,-81</points>
<connection>
<GID>336</GID>
<name>IN_1</name></connection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70,-64,81,-64</points>
<connection>
<GID>305</GID>
<name>OUT</name></connection>
<intersection>81 0</intersection></hsegment></shape></wire>
<wire>
<ID>209</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82,-67,82,-60</points>
<intersection>-67 1</intersection>
<intersection>-60 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82,-67,104,-67</points>
<connection>
<GID>335</GID>
<name>IN_1</name></connection>
<intersection>82 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70,-60,82,-60</points>
<connection>
<GID>304</GID>
<name>OUT</name></connection>
<intersection>82 0</intersection></hsegment></shape></wire>
<wire>
<ID>210</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82,-56,82,-53</points>
<intersection>-56 2</intersection>
<intersection>-53 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82,-53,104,-53</points>
<connection>
<GID>334</GID>
<name>IN_1</name></connection>
<intersection>82 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70,-56,82,-56</points>
<connection>
<GID>303</GID>
<name>OUT</name></connection>
<intersection>82 0</intersection></hsegment></shape></wire>
<wire>
<ID>211</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82,-52,82,-39</points>
<intersection>-52 2</intersection>
<intersection>-39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82,-39,104,-39</points>
<connection>
<GID>333</GID>
<name>IN_1</name></connection>
<intersection>82 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70,-52,82,-52</points>
<connection>
<GID>302</GID>
<name>OUT</name></connection>
<intersection>82 0</intersection></hsegment></shape></wire>
<wire>
<ID>212</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,-48,81,-25</points>
<intersection>-48 2</intersection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>81,-25,104,-25</points>
<connection>
<GID>332</GID>
<name>IN_1</name></connection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70,-48,81,-48</points>
<connection>
<GID>301</GID>
<name>OUT</name></connection>
<intersection>81 0</intersection></hsegment></shape></wire>
<wire>
<ID>213</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78,-27,78,-14</points>
<intersection>-27 1</intersection>
<intersection>-14 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>78,-27,104,-27</points>
<connection>
<GID>332</GID>
<name>IN_0</name></connection>
<intersection>78 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70,-14,78,-14</points>
<connection>
<GID>292</GID>
<name>OUT</name></connection>
<intersection>78 0</intersection></hsegment></shape></wire>
<wire>
<ID>214</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71,-125,71,-42</points>
<intersection>-125 1</intersection>
<intersection>-42 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>71,-125,104,-125</points>
<connection>
<GID>339</GID>
<name>IN_0</name></connection>
<intersection>71 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70,-42,71,-42</points>
<connection>
<GID>299</GID>
<name>OUT</name></connection>
<intersection>71 0</intersection></hsegment></shape></wire>
<wire>
<ID>215</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-111,72,-38</points>
<intersection>-111 1</intersection>
<intersection>-38 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72,-111,104,-111</points>
<connection>
<GID>338</GID>
<name>IN_0</name></connection>
<intersection>72 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70,-38,72,-38</points>
<connection>
<GID>298</GID>
<name>OUT</name></connection>
<intersection>72 0</intersection></hsegment></shape></wire>
<wire>
<ID>216</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-97,73,-34</points>
<intersection>-97 1</intersection>
<intersection>-34 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73,-97,104,-97</points>
<connection>
<GID>337</GID>
<name>IN_0</name></connection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70,-34,73,-34</points>
<connection>
<GID>297</GID>
<name>OUT</name></connection>
<intersection>73 0</intersection></hsegment></shape></wire>
<wire>
<ID>217</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74,-83,74,-30</points>
<intersection>-83 1</intersection>
<intersection>-30 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74,-83,104,-83</points>
<connection>
<GID>336</GID>
<name>IN_0</name></connection>
<intersection>74 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70,-30,74,-30</points>
<connection>
<GID>296</GID>
<name>OUT</name></connection>
<intersection>74 0</intersection></hsegment></shape></wire>
<wire>
<ID>218</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-69,75,-26</points>
<intersection>-69 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75,-69,104,-69</points>
<connection>
<GID>335</GID>
<name>IN_0</name></connection>
<intersection>75 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70,-26,75,-26</points>
<connection>
<GID>295</GID>
<name>OUT</name></connection>
<intersection>75 0</intersection></hsegment></shape></wire>
<wire>
<ID>220</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-55,76,-22</points>
<intersection>-55 1</intersection>
<intersection>-22 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76,-55,104,-55</points>
<connection>
<GID>334</GID>
<name>IN_0</name></connection>
<intersection>76 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70,-22,76,-22</points>
<connection>
<GID>294</GID>
<name>OUT</name></connection>
<intersection>76 0</intersection></hsegment></shape></wire>
<wire>
<ID>221</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77,-41,77,-18</points>
<intersection>-41 1</intersection>
<intersection>-18 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77,-41,104,-41</points>
<connection>
<GID>333</GID>
<name>IN_0</name></connection>
<intersection>77 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70,-18,77,-18</points>
<connection>
<GID>293</GID>
<name>OUT</name></connection>
<intersection>77 0</intersection></hsegment></shape></wire>
<wire>
<ID>222</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117,-117,117,-9</points>
<intersection>-117 3</intersection>
<intersection>-103 4</intersection>
<intersection>-89 7</intersection>
<intersection>-75 8</intersection>
<intersection>-61 9</intersection>
<intersection>-47 10</intersection>
<intersection>-33 11</intersection>
<intersection>-19 12</intersection>
<intersection>-9 5</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>108,-117,117,-117</points>
<connection>
<GID>339</GID>
<name>SEL_0</name></connection>
<intersection>117 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>108,-103,117,-103</points>
<connection>
<GID>338</GID>
<name>SEL_0</name></connection>
<intersection>117 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>117,-9,118,-9</points>
<intersection>117 0</intersection>
<intersection>118 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>118,-9,118,-7</points>
<connection>
<GID>259</GID>
<name>OUT_0</name></connection>
<intersection>-9 5</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>108,-89,117,-89</points>
<connection>
<GID>337</GID>
<name>SEL_0</name></connection>
<intersection>117 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>108,-75,117,-75</points>
<connection>
<GID>336</GID>
<name>SEL_0</name></connection>
<intersection>117 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>108,-61,117,-61</points>
<connection>
<GID>335</GID>
<name>SEL_0</name></connection>
<intersection>117 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>108,-47,117,-47</points>
<connection>
<GID>334</GID>
<name>SEL_0</name></connection>
<intersection>117 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>108,-33,117,-33</points>
<connection>
<GID>333</GID>
<name>SEL_0</name></connection>
<intersection>117 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>108,-19,117,-19</points>
<connection>
<GID>332</GID>
<name>SEL_0</name></connection>
<intersection>117 0</intersection></hsegment></shape></wire>
<wire>
<ID>223</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116,-116,116,-9</points>
<intersection>-116 3</intersection>
<intersection>-102 7</intersection>
<intersection>-88 9</intersection>
<intersection>-74 11</intersection>
<intersection>-60 13</intersection>
<intersection>-46 15</intersection>
<intersection>-32 17</intersection>
<intersection>-18 19</intersection>
<intersection>-9 5</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>107,-116,116,-116</points>
<intersection>107 21</intersection>
<intersection>116 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>115,-9,116,-9</points>
<intersection>115 6</intersection>
<intersection>116 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>115,-9,115,-7</points>
<connection>
<GID>258</GID>
<name>OUT_0</name></connection>
<intersection>-9 5</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>107,-102,116,-102</points>
<intersection>107 8</intersection>
<intersection>116 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>107,-103,107,-102</points>
<connection>
<GID>338</GID>
<name>SEL_1</name></connection>
<intersection>-102 7</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>107,-88,116,-88</points>
<intersection>107 10</intersection>
<intersection>116 0</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>107,-89,107,-88</points>
<connection>
<GID>337</GID>
<name>SEL_1</name></connection>
<intersection>-88 9</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>107,-74,116,-74</points>
<intersection>107 12</intersection>
<intersection>116 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>107,-75,107,-74</points>
<connection>
<GID>336</GID>
<name>SEL_1</name></connection>
<intersection>-74 11</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>107,-60,116,-60</points>
<intersection>107 14</intersection>
<intersection>116 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>107,-61,107,-60</points>
<connection>
<GID>335</GID>
<name>SEL_1</name></connection>
<intersection>-60 13</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>107,-46,116,-46</points>
<intersection>107 16</intersection>
<intersection>116 0</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>107,-47,107,-46</points>
<connection>
<GID>334</GID>
<name>SEL_1</name></connection>
<intersection>-46 15</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>107,-32,116,-32</points>
<intersection>107 18</intersection>
<intersection>116 0</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>107,-33,107,-32</points>
<connection>
<GID>333</GID>
<name>SEL_1</name></connection>
<intersection>-32 17</intersection></vsegment>
<hsegment>
<ID>19</ID>
<points>107,-18,116,-18</points>
<intersection>107 20</intersection>
<intersection>116 0</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>107,-19,107,-18</points>
<connection>
<GID>332</GID>
<name>SEL_1</name></connection>
<intersection>-18 19</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>107,-117,107,-116</points>
<connection>
<GID>339</GID>
<name>SEL_1</name></connection>
<intersection>-116 3</intersection></vsegment></shape></wire>
<wire>
<ID>224</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127,-59,127,-24</points>
<intersection>-59 1</intersection>
<intersection>-24 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127,-59,129,-59</points>
<connection>
<GID>234</GID>
<name>N_in0</name></connection>
<intersection>127 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>110,-24,127,-24</points>
<connection>
<GID>332</GID>
<name>OUT</name></connection>
<intersection>127 0</intersection></hsegment></shape></wire>
<wire>
<ID>225</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,-63,125,-38</points>
<intersection>-63 1</intersection>
<intersection>-38 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>125,-63,129,-63</points>
<connection>
<GID>235</GID>
<name>N_in0</name></connection>
<intersection>125 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>110,-38,125,-38</points>
<connection>
<GID>333</GID>
<name>OUT</name></connection>
<intersection>125 0</intersection></hsegment></shape></wire>
<wire>
<ID>226</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123,-67,123,-52</points>
<intersection>-67 1</intersection>
<intersection>-52 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123,-67,129,-67</points>
<connection>
<GID>236</GID>
<name>N_in0</name></connection>
<intersection>123 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>110,-52,123,-52</points>
<connection>
<GID>334</GID>
<name>OUT</name></connection>
<intersection>123 0</intersection></hsegment></shape></wire>
<wire>
<ID>227</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121,-71,121,-66</points>
<intersection>-71 1</intersection>
<intersection>-66 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121,-71,129,-71</points>
<connection>
<GID>237</GID>
<name>N_in0</name></connection>
<intersection>121 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>110,-66,121,-66</points>
<connection>
<GID>335</GID>
<name>OUT</name></connection>
<intersection>121 0</intersection></hsegment></shape></wire>
<wire>
<ID>228</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121,-80,121,-75</points>
<intersection>-80 2</intersection>
<intersection>-75 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121,-75,129,-75</points>
<connection>
<GID>243</GID>
<name>N_in0</name></connection>
<intersection>121 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>110,-80,121,-80</points>
<connection>
<GID>336</GID>
<name>OUT</name></connection>
<intersection>121 0</intersection></hsegment></shape></wire>
<wire>
<ID>229</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123,-94,123,-79</points>
<intersection>-94 2</intersection>
<intersection>-79 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123,-79,129,-79</points>
<connection>
<GID>244</GID>
<name>N_in0</name></connection>
<intersection>123 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>110,-94,123,-94</points>
<connection>
<GID>337</GID>
<name>OUT</name></connection>
<intersection>123 0</intersection></hsegment></shape></wire>
<wire>
<ID>230</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,-108,125,-83</points>
<intersection>-108 2</intersection>
<intersection>-83 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>125,-83,129,-83</points>
<connection>
<GID>245</GID>
<name>N_in0</name></connection>
<intersection>125 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>110,-108,125,-108</points>
<connection>
<GID>338</GID>
<name>OUT</name></connection>
<intersection>125 0</intersection></hsegment></shape></wire>
<wire>
<ID>231</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127,-122,127,-87</points>
<intersection>-122 2</intersection>
<intersection>-87 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127,-87,129,-87</points>
<connection>
<GID>246</GID>
<name>N_in0</name></connection>
<intersection>127 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>110,-122,127,-122</points>
<connection>
<GID>339</GID>
<name>OUT</name></connection>
<intersection>127 0</intersection></hsegment></shape></wire>
<wire>
<ID>235</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-81,40,-7</points>
<connection>
<GID>205</GID>
<name>OUT_0</name></connection>
<intersection>-81 1</intersection>
<intersection>-47 2</intersection>
<intersection>-13 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,-81,64.5,-81</points>
<connection>
<GID>310</GID>
<name>IN_0</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>40,-47,64,-47</points>
<connection>
<GID>301</GID>
<name>IN_0</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>40,-13,64,-13</points>
<connection>
<GID>292</GID>
<name>IN_0</name></connection>
<intersection>40 0</intersection></hsegment></shape></wire>
<wire>
<ID>236</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10,-116,10,-7</points>
<connection>
<GID>247</GID>
<name>OUT_0</name></connection>
<intersection>-116 7</intersection>
<intersection>-83 1</intersection>
<intersection>-49 3</intersection>
<intersection>-15 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10,-83,64.5,-83</points>
<connection>
<GID>310</GID>
<name>IN_1</name></connection>
<intersection>10 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>10,-49,64,-49</points>
<connection>
<GID>301</GID>
<name>IN_1</name></connection>
<intersection>10 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>10,-15,64,-15</points>
<connection>
<GID>292</GID>
<name>IN_1</name></connection>
<intersection>10 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>10,-116,65,-116</points>
<connection>
<GID>323</GID>
<name>IN_0</name></connection>
<intersection>10 0</intersection></hsegment></shape></wire>
<wire>
<ID>237</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43,-85,43,-7</points>
<connection>
<GID>206</GID>
<name>OUT_0</name></connection>
<intersection>-85 1</intersection>
<intersection>-51 2</intersection>
<intersection>-17 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43,-85,64.5,-85</points>
<connection>
<GID>311</GID>
<name>IN_0</name></connection>
<intersection>43 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43,-51,64,-51</points>
<connection>
<GID>302</GID>
<name>IN_0</name></connection>
<intersection>43 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>43,-17,64,-17</points>
<connection>
<GID>293</GID>
<name>IN_0</name></connection>
<intersection>43 0</intersection></hsegment></shape></wire>
<wire>
<ID>238</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-119,13,-7</points>
<connection>
<GID>248</GID>
<name>OUT_0</name></connection>
<intersection>-119 7</intersection>
<intersection>-87 1</intersection>
<intersection>-53 3</intersection>
<intersection>-19 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13,-87,64.5,-87</points>
<connection>
<GID>311</GID>
<name>IN_1</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>13,-53,64,-53</points>
<connection>
<GID>302</GID>
<name>IN_1</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>13,-19,64,-19</points>
<connection>
<GID>293</GID>
<name>IN_1</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>13,-119,65,-119</points>
<connection>
<GID>324</GID>
<name>IN_0</name></connection>
<intersection>13 0</intersection></hsegment></shape></wire>
<wire>
<ID>239</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-89,46,-7</points>
<connection>
<GID>207</GID>
<name>OUT_0</name></connection>
<intersection>-89 1</intersection>
<intersection>-55 2</intersection>
<intersection>-21 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-89,64.5,-89</points>
<connection>
<GID>312</GID>
<name>IN_0</name></connection>
<intersection>46 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>46,-55,64,-55</points>
<connection>
<GID>303</GID>
<name>IN_0</name></connection>
<intersection>46 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>46,-21,64,-21</points>
<connection>
<GID>294</GID>
<name>IN_0</name></connection>
<intersection>46 0</intersection></hsegment></shape></wire>
<wire>
<ID>240</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16,-122,16,-7</points>
<connection>
<GID>249</GID>
<name>OUT_0</name></connection>
<intersection>-122 7</intersection>
<intersection>-91 1</intersection>
<intersection>-57 3</intersection>
<intersection>-23 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16,-91,64.5,-91</points>
<connection>
<GID>312</GID>
<name>IN_1</name></connection>
<intersection>16 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>16,-57,64,-57</points>
<connection>
<GID>303</GID>
<name>IN_1</name></connection>
<intersection>16 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>16,-23,64,-23</points>
<connection>
<GID>294</GID>
<name>IN_1</name></connection>
<intersection>16 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>16,-122,65,-122</points>
<connection>
<GID>325</GID>
<name>IN_0</name></connection>
<intersection>16 0</intersection></hsegment></shape></wire>
<wire>
<ID>241</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49,-93,49,-7</points>
<connection>
<GID>208</GID>
<name>OUT_0</name></connection>
<intersection>-93 1</intersection>
<intersection>-59 2</intersection>
<intersection>-25 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49,-93,64.5,-93</points>
<connection>
<GID>313</GID>
<name>IN_0</name></connection>
<intersection>49 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49,-59,64,-59</points>
<connection>
<GID>304</GID>
<name>IN_0</name></connection>
<intersection>49 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>49,-25,64,-25</points>
<connection>
<GID>295</GID>
<name>IN_0</name></connection>
<intersection>49 0</intersection></hsegment></shape></wire>
<wire>
<ID>242</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,-125,19,-7</points>
<connection>
<GID>250</GID>
<name>OUT_0</name></connection>
<intersection>-125 7</intersection>
<intersection>-95 1</intersection>
<intersection>-61 3</intersection>
<intersection>-27 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19,-95,64.5,-95</points>
<connection>
<GID>313</GID>
<name>IN_1</name></connection>
<intersection>19 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>19,-61,64,-61</points>
<connection>
<GID>304</GID>
<name>IN_1</name></connection>
<intersection>19 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>19,-27,64,-27</points>
<connection>
<GID>295</GID>
<name>IN_1</name></connection>
<intersection>19 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>19,-125,65,-125</points>
<connection>
<GID>326</GID>
<name>IN_0</name></connection>
<intersection>19 0</intersection></hsegment></shape></wire>
<wire>
<ID>243</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-97,52,-7</points>
<connection>
<GID>209</GID>
<name>OUT_0</name></connection>
<intersection>-97 1</intersection>
<intersection>-63 2</intersection>
<intersection>-29 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52,-97,64.5,-97</points>
<connection>
<GID>314</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>52,-63,64,-63</points>
<connection>
<GID>305</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>52,-29,64,-29</points>
<connection>
<GID>296</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>244</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-128,21.5,-7</points>
<connection>
<GID>251</GID>
<name>OUT_0</name></connection>
<intersection>-128 7</intersection>
<intersection>-99 1</intersection>
<intersection>-65 3</intersection>
<intersection>-31 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21.5,-99,64.5,-99</points>
<connection>
<GID>314</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>21.5,-65,64,-65</points>
<connection>
<GID>305</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>21.5,-31,64,-31</points>
<connection>
<GID>296</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>21.5,-128,65,-128</points>
<connection>
<GID>327</GID>
<name>IN_0</name></connection>
<intersection>21.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>245</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55,-101,55,-7</points>
<connection>
<GID>210</GID>
<name>OUT_0</name></connection>
<intersection>-101 1</intersection>
<intersection>-67 2</intersection>
<intersection>-33 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55,-101,64.5,-101</points>
<connection>
<GID>315</GID>
<name>IN_0</name></connection>
<intersection>55 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>55,-67,64,-67</points>
<connection>
<GID>306</GID>
<name>IN_0</name></connection>
<intersection>55 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>55,-33,64,-33</points>
<connection>
<GID>297</GID>
<name>IN_0</name></connection>
<intersection>55 0</intersection></hsegment></shape></wire>
<wire>
<ID>246</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-131,25,-7</points>
<connection>
<GID>252</GID>
<name>OUT_0</name></connection>
<intersection>-131 7</intersection>
<intersection>-103 1</intersection>
<intersection>-69 3</intersection>
<intersection>-35 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-103,64.5,-103</points>
<connection>
<GID>315</GID>
<name>IN_1</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>25,-69,64,-69</points>
<connection>
<GID>306</GID>
<name>IN_1</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>25,-35,64,-35</points>
<connection>
<GID>297</GID>
<name>IN_1</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>25,-131,65,-131</points>
<connection>
<GID>328</GID>
<name>IN_0</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>247</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58,-105,58,-7</points>
<connection>
<GID>211</GID>
<name>OUT_0</name></connection>
<intersection>-105 1</intersection>
<intersection>-71 2</intersection>
<intersection>-37 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58,-105,64.5,-105</points>
<connection>
<GID>316</GID>
<name>IN_0</name></connection>
<intersection>58 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>58,-71,64,-71</points>
<connection>
<GID>307</GID>
<name>IN_0</name></connection>
<intersection>58 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>58,-37,64,-37</points>
<connection>
<GID>298</GID>
<name>IN_0</name></connection>
<intersection>58 0</intersection></hsegment></shape></wire>
<wire>
<ID>248</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-134,28,-7</points>
<connection>
<GID>253</GID>
<name>OUT_0</name></connection>
<intersection>-134 7</intersection>
<intersection>-107 1</intersection>
<intersection>-73 3</intersection>
<intersection>-39 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-107,64.5,-107</points>
<connection>
<GID>316</GID>
<name>IN_1</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>28,-73,64,-73</points>
<connection>
<GID>307</GID>
<name>IN_1</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>28,-39,64,-39</points>
<connection>
<GID>298</GID>
<name>IN_1</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>28,-134,65,-134</points>
<connection>
<GID>329</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>249</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-109,61,-7</points>
<connection>
<GID>212</GID>
<name>OUT_0</name></connection>
<intersection>-109 1</intersection>
<intersection>-75 2</intersection>
<intersection>-41 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61,-109,64.5,-109</points>
<connection>
<GID>317</GID>
<name>IN_0</name></connection>
<intersection>61 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>61,-75,64,-75</points>
<connection>
<GID>308</GID>
<name>IN_0</name></connection>
<intersection>61 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>61,-41,64,-41</points>
<connection>
<GID>299</GID>
<name>IN_0</name></connection>
<intersection>61 0</intersection></hsegment></shape></wire>
<wire>
<ID>250</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-137,31,-7</points>
<connection>
<GID>254</GID>
<name>OUT_0</name></connection>
<intersection>-137 5</intersection>
<intersection>-111 1</intersection>
<intersection>-77 2</intersection>
<intersection>-43 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-111,64.5,-111</points>
<connection>
<GID>317</GID>
<name>IN_1</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31,-77,64,-77</points>
<connection>
<GID>308</GID>
<name>IN_1</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>31,-43,64,-43</points>
<connection>
<GID>299</GID>
<name>IN_1</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>31,-137,65,-137</points>
<connection>
<GID>330</GID>
<name>IN_0</name></connection>
<intersection>31 0</intersection></hsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93,-116,93,-21</points>
<intersection>-116 2</intersection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>93,-21,104,-21</points>
<connection>
<GID>332</GID>
<name>IN_3</name></connection>
<intersection>93 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69,-116,93,-116</points>
<connection>
<GID>323</GID>
<name>OUT_0</name></connection>
<intersection>93 0</intersection></hsegment></shape></wire>
<wire>
<ID>190</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>94,-119,94,-35</points>
<intersection>-119 2</intersection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>94,-35,104,-35</points>
<connection>
<GID>333</GID>
<name>IN_3</name></connection>
<intersection>94 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69,-119,94,-119</points>
<connection>
<GID>324</GID>
<name>OUT_0</name></connection>
<intersection>94 0</intersection></hsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95,-122,95,-49</points>
<intersection>-122 2</intersection>
<intersection>-49 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95,-49,104,-49</points>
<connection>
<GID>334</GID>
<name>IN_3</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69,-122,95,-122</points>
<connection>
<GID>325</GID>
<name>OUT_0</name></connection>
<intersection>95 0</intersection></hsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96,-125,96,-63</points>
<intersection>-125 2</intersection>
<intersection>-63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>96,-63,104,-63</points>
<connection>
<GID>335</GID>
<name>IN_3</name></connection>
<intersection>96 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69,-125,96,-125</points>
<connection>
<GID>326</GID>
<name>OUT_0</name></connection>
<intersection>96 0</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>-22.0087,-45.4589,458.684,-293.375</PageViewport>
<gate>
<ID>389</ID>
<type>AA_LABEL</type>
<position>302,-147.5</position>
<gparam>LABEL_TEXT G0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>390</ID>
<type>GA_LED</type>
<position>299.5,-120</position>
<input>
<ID>N_in0</ID>181 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1</ID>
<type>AA_TOGGLE</type>
<position>225.5,-66</position>
<output>
<ID>OUT_0</ID>256 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>391</ID>
<type>GA_LED</type>
<position>299.5,-124</position>
<input>
<ID>N_in0</ID>182 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>225.5,-63.5</position>
<gparam>LABEL_TEXT S3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>392</ID>
<type>GA_LED</type>
<position>299.5,-128</position>
<input>
<ID>N_in0</ID>183 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3</ID>
<type>AA_TOGGLE</type>
<position>148,-66</position>
<output>
<ID>OUT_0</ID>61 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>393</ID>
<type>GA_LED</type>
<position>299.5,-132</position>
<input>
<ID>N_in0</ID>184 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>151,-66</position>
<output>
<ID>OUT_0</ID>63 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>394</ID>
<type>AA_LABEL</type>
<position>302,-120</position>
<gparam>LABEL_TEXT G7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>5</ID>
<type>AA_TOGGLE</type>
<position>154,-66</position>
<output>
<ID>OUT_0</ID>257 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>395</ID>
<type>AA_LABEL</type>
<position>302,-124</position>
<gparam>LABEL_TEXT G6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>157,-66</position>
<output>
<ID>OUT_0</ID>110 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>396</ID>
<type>AA_LABEL</type>
<position>302,-128</position>
<gparam>LABEL_TEXT G5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7</ID>
<type>AA_TOGGLE</type>
<position>160,-66</position>
<output>
<ID>OUT_0</ID>112 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>397</ID>
<type>AA_LABEL</type>
<position>302,-132</position>
<gparam>LABEL_TEXT G4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>163,-66</position>
<output>
<ID>OUT_0</ID>114 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>398</ID>
<type>GA_LED</type>
<position>299.5,-136</position>
<input>
<ID>N_in0</ID>185 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>9</ID>
<type>AA_TOGGLE</type>
<position>166,-66</position>
<output>
<ID>OUT_0</ID>116 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>399</ID>
<type>GA_LED</type>
<position>299.5,-140</position>
<input>
<ID>N_in0</ID>186 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>169,-66</position>
<output>
<ID>OUT_0</ID>118 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>400</ID>
<type>GA_LED</type>
<position>299.5,-144</position>
<input>
<ID>N_in0</ID>187 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>AA_LABEL</type>
<position>118,-63.5</position>
<gparam>LABEL_TEXT X7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>401</ID>
<type>GA_LED</type>
<position>299.5,-148</position>
<input>
<ID>N_in0</ID>188 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AA_LABEL</type>
<position>121,-63.5</position>
<gparam>LABEL_TEXT X6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>13</ID>
<type>AA_LABEL</type>
<position>124,-63.5</position>
<gparam>LABEL_TEXT X5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>403</ID>
<type>AA_LABEL</type>
<position>299.5,-111.5</position>
<gparam>LABEL_TEXT Cout</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>AA_LABEL</type>
<position>127,-63.5</position>
<gparam>LABEL_TEXT X4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>404</ID>
<type>GA_LED</type>
<position>299.5,-114</position>
<input>
<ID>N_in1</ID>268 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>AA_LABEL</type>
<position>130,-63.5</position>
<gparam>LABEL_TEXT X3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>AA_LABEL</type>
<position>133,-63.5</position>
<gparam>LABEL_TEXT X2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>17</ID>
<type>AA_LABEL</type>
<position>136,-63.5</position>
<gparam>LABEL_TEXT X1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>408</ID>
<type>AA_LABEL</type>
<position>203,-47</position>
<gparam>LABEL_TEXT Unidade Logica e Aritmetica</gparam>
<gparam>TEXT_HEIGHT 5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>AA_LABEL</type>
<position>139,-63.5</position>
<gparam>LABEL_TEXT X0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>21</ID>
<type>AA_LABEL</type>
<position>148,-63.5</position>
<gparam>LABEL_TEXT Y7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>23</ID>
<type>AA_LABEL</type>
<position>151,-63.5</position>
<gparam>LABEL_TEXT Y6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>25</ID>
<type>AA_LABEL</type>
<position>154,-63.5</position>
<gparam>LABEL_TEXT Y5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>27</ID>
<type>AA_LABEL</type>
<position>157,-63.5</position>
<gparam>LABEL_TEXT Y4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>AA_LABEL</type>
<position>160,-63.5</position>
<gparam>LABEL_TEXT Y3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>AA_LABEL</type>
<position>163,-63.5</position>
<gparam>LABEL_TEXT Y2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>33</ID>
<type>AA_LABEL</type>
<position>166,-63.5</position>
<gparam>LABEL_TEXT Y1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>50</ID>
<type>AA_LABEL</type>
<position>169,-63.5</position>
<gparam>LABEL_TEXT Y0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>71</ID>
<type>AA_TOGGLE</type>
<position>118,-66</position>
<output>
<ID>OUT_0</ID>62 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>72</ID>
<type>AA_TOGGLE</type>
<position>121,-66</position>
<output>
<ID>OUT_0</ID>81 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>73</ID>
<type>AA_TOGGLE</type>
<position>124,-66</position>
<output>
<ID>OUT_0</ID>109 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>74</ID>
<type>AA_TOGGLE</type>
<position>127,-66</position>
<output>
<ID>OUT_0</ID>111 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>75</ID>
<type>AA_TOGGLE</type>
<position>130,-66</position>
<output>
<ID>OUT_0</ID>113 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>76</ID>
<type>AA_TOGGLE</type>
<position>133,-66</position>
<output>
<ID>OUT_0</ID>115 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>77</ID>
<type>AA_TOGGLE</type>
<position>136,-66</position>
<output>
<ID>OUT_0</ID>117 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>78</ID>
<type>AA_TOGGLE</type>
<position>139,-66</position>
<output>
<ID>OUT_0</ID>119 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>79</ID>
<type>AA_TOGGLE</type>
<position>228.5,-66</position>
<output>
<ID>OUT_0</ID>259 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>80</ID>
<type>AA_TOGGLE</type>
<position>231.5,-66</position>
<output>
<ID>OUT_0</ID>258 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>81</ID>
<type>AA_TOGGLE</type>
<position>234.5,-66</position>
<output>
<ID>OUT_0</ID>41 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>83</ID>
<type>AA_LABEL</type>
<position>228.5,-63.5</position>
<gparam>LABEL_TEXT S2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>85</ID>
<type>AA_LABEL</type>
<position>231.5,-63.5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>87</ID>
<type>AA_LABEL</type>
<position>234.5,-63.5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>89</ID>
<type>AA_AND2</type>
<position>175,-75</position>
<input>
<ID>IN_0</ID>61 </input>
<input>
<ID>IN_1</ID>62 </input>
<output>
<ID>OUT</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>91</ID>
<type>AA_AND2</type>
<position>175,-79</position>
<input>
<ID>IN_0</ID>63 </input>
<input>
<ID>IN_1</ID>81 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>109</ID>
<type>AA_AND2</type>
<position>175,-83</position>
<input>
<ID>IN_0</ID>257 </input>
<input>
<ID>IN_1</ID>109 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>110</ID>
<type>AA_AND2</type>
<position>175,-87</position>
<input>
<ID>IN_0</ID>110 </input>
<input>
<ID>IN_1</ID>111 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>111</ID>
<type>AA_AND2</type>
<position>175,-91</position>
<input>
<ID>IN_0</ID>112 </input>
<input>
<ID>IN_1</ID>113 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>112</ID>
<type>AA_AND2</type>
<position>175,-95</position>
<input>
<ID>IN_0</ID>114 </input>
<input>
<ID>IN_1</ID>115 </input>
<output>
<ID>OUT</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>113</ID>
<type>AA_AND2</type>
<position>175,-99</position>
<input>
<ID>IN_0</ID>116 </input>
<input>
<ID>IN_1</ID>117 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>114</ID>
<type>AA_AND2</type>
<position>175,-103</position>
<input>
<ID>IN_0</ID>118 </input>
<input>
<ID>IN_1</ID>119 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>115</ID>
<type>AE_OR2</type>
<position>175,-109</position>
<input>
<ID>IN_0</ID>61 </input>
<input>
<ID>IN_1</ID>62 </input>
<output>
<ID>OUT</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>116</ID>
<type>AE_OR2</type>
<position>175,-113</position>
<input>
<ID>IN_0</ID>63 </input>
<input>
<ID>IN_1</ID>81 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>117</ID>
<type>AE_OR2</type>
<position>175,-117</position>
<input>
<ID>IN_0</ID>257 </input>
<input>
<ID>IN_1</ID>109 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>118</ID>
<type>AE_OR2</type>
<position>175,-121</position>
<input>
<ID>IN_0</ID>110 </input>
<input>
<ID>IN_1</ID>111 </input>
<output>
<ID>OUT</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>119</ID>
<type>AE_OR2</type>
<position>175,-125</position>
<input>
<ID>IN_0</ID>112 </input>
<input>
<ID>IN_1</ID>113 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>120</ID>
<type>AE_OR2</type>
<position>175,-129</position>
<input>
<ID>IN_0</ID>114 </input>
<input>
<ID>IN_1</ID>115 </input>
<output>
<ID>OUT</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>121</ID>
<type>AE_OR2</type>
<position>175,-133</position>
<input>
<ID>IN_0</ID>116 </input>
<input>
<ID>IN_1</ID>117 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>122</ID>
<type>AE_OR2</type>
<position>175,-137</position>
<input>
<ID>IN_0</ID>118 </input>
<input>
<ID>IN_1</ID>119 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>512</ID>
<type>AA_LABEL</type>
<position>128.5,-60</position>
<gparam>LABEL_TEXT Entradas (X)</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>123</ID>
<type>AI_XOR2</type>
<position>175.5,-143</position>
<input>
<ID>IN_0</ID>61 </input>
<input>
<ID>IN_1</ID>62 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>513</ID>
<type>AA_LABEL</type>
<position>158.5,-60</position>
<gparam>LABEL_TEXT Entradas (Y)</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>124</ID>
<type>AI_XOR2</type>
<position>175.5,-147</position>
<input>
<ID>IN_0</ID>63 </input>
<input>
<ID>IN_1</ID>81 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>514</ID>
<type>AA_LABEL</type>
<position>230,-60</position>
<gparam>LABEL_TEXT Seletores (S)</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>125</ID>
<type>AI_XOR2</type>
<position>175.5,-151</position>
<input>
<ID>IN_0</ID>257 </input>
<input>
<ID>IN_1</ID>109 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>515</ID>
<type>AA_LABEL</type>
<position>315,-130.5</position>
<gparam>LABEL_TEXT Saidas (G)</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>126</ID>
<type>AI_XOR2</type>
<position>175.5,-155</position>
<input>
<ID>IN_0</ID>110 </input>
<input>
<ID>IN_1</ID>111 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>516</ID>
<type>AA_LABEL</type>
<position>175,-72</position>
<gparam>LABEL_TEXT 74HC08</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>127</ID>
<type>AI_XOR2</type>
<position>175.5,-159</position>
<input>
<ID>IN_0</ID>112 </input>
<input>
<ID>IN_1</ID>113 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>517</ID>
<type>AA_LABEL</type>
<position>175,-106</position>
<gparam>LABEL_TEXT 74HC32</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>128</ID>
<type>AI_XOR2</type>
<position>175.5,-163</position>
<input>
<ID>IN_0</ID>114 </input>
<input>
<ID>IN_1</ID>115 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>518</ID>
<type>AA_LABEL</type>
<position>175,-140</position>
<gparam>LABEL_TEXT 74HC86</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>129</ID>
<type>AI_XOR2</type>
<position>175.5,-167</position>
<input>
<ID>IN_0</ID>116 </input>
<input>
<ID>IN_1</ID>117 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>519</ID>
<type>AA_LABEL</type>
<position>175,-175</position>
<gparam>LABEL_TEXT 74HC04</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>130</ID>
<type>AI_XOR2</type>
<position>175.5,-171</position>
<input>
<ID>IN_0</ID>118 </input>
<input>
<ID>IN_1</ID>119 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>520</ID>
<type>AA_LABEL</type>
<position>170.5,-75</position>
<gparam>LABEL_TEXT U1a</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>131</ID>
<type>AE_SMALL_INVERTER</type>
<position>175,-177</position>
<input>
<ID>IN_0</ID>62 </input>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>521</ID>
<type>AA_LABEL</type>
<position>170.5,-79</position>
<gparam>LABEL_TEXT U1b</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>132</ID>
<type>AE_SMALL_INVERTER</type>
<position>175,-180</position>
<input>
<ID>IN_0</ID>81 </input>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>522</ID>
<type>AA_LABEL</type>
<position>170.5,-83</position>
<gparam>LABEL_TEXT U1c</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>133</ID>
<type>AE_SMALL_INVERTER</type>
<position>175,-183</position>
<input>
<ID>IN_0</ID>109 </input>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>523</ID>
<type>AA_LABEL</type>
<position>170.5,-87</position>
<gparam>LABEL_TEXT U1d</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>134</ID>
<type>AE_SMALL_INVERTER</type>
<position>175,-186</position>
<input>
<ID>IN_0</ID>111 </input>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>524</ID>
<type>AA_LABEL</type>
<position>170.5,-91</position>
<gparam>LABEL_TEXT U1e</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>135</ID>
<type>AE_SMALL_INVERTER</type>
<position>175,-189</position>
<input>
<ID>IN_0</ID>113 </input>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>525</ID>
<type>AA_LABEL</type>
<position>170.5,-95</position>
<gparam>LABEL_TEXT U1f</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>136</ID>
<type>AE_SMALL_INVERTER</type>
<position>175,-192</position>
<input>
<ID>IN_0</ID>115 </input>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>526</ID>
<type>AA_LABEL</type>
<position>170.5,-99</position>
<gparam>LABEL_TEXT U1g</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>137</ID>
<type>AE_SMALL_INVERTER</type>
<position>175,-195</position>
<input>
<ID>IN_0</ID>117 </input>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>527</ID>
<type>AA_LABEL</type>
<position>170.5,-103</position>
<gparam>LABEL_TEXT U1h</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>528</ID>
<type>AA_LABEL</type>
<position>170.5,-109</position>
<gparam>LABEL_TEXT U2a</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>529</ID>
<type>AA_LABEL</type>
<position>170.5,-113</position>
<gparam>LABEL_TEXT U2b</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>140</ID>
<type>AE_SMALL_INVERTER</type>
<position>175,-198</position>
<input>
<ID>IN_0</ID>119 </input>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>530</ID>
<type>AA_LABEL</type>
<position>170.5,-117</position>
<gparam>LABEL_TEXT U2c</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>141</ID>
<type>AE_MUX_4x1</type>
<position>217,-85</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>24 </input>
<input>
<ID>IN_2</ID>9 </input>
<input>
<ID>IN_3</ID>1 </input>
<output>
<ID>OUT</ID>219 </output>
<input>
<ID>SEL_0</ID>41 </input>
<input>
<ID>SEL_1</ID>258 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>531</ID>
<type>AA_LABEL</type>
<position>170.5,-121</position>
<gparam>LABEL_TEXT U2d</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>142</ID>
<type>AE_MUX_4x1</type>
<position>217,-99</position>
<input>
<ID>IN_0</ID>40 </input>
<input>
<ID>IN_1</ID>23 </input>
<input>
<ID>IN_2</ID>16 </input>
<input>
<ID>IN_3</ID>2 </input>
<output>
<ID>OUT</ID>255 </output>
<input>
<ID>SEL_0</ID>41 </input>
<input>
<ID>SEL_1</ID>258 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>532</ID>
<type>AA_LABEL</type>
<position>170.5,-125</position>
<gparam>LABEL_TEXT U2e</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>143</ID>
<type>AE_MUX_4x1</type>
<position>217,-113</position>
<input>
<ID>IN_0</ID>39 </input>
<input>
<ID>IN_1</ID>22 </input>
<input>
<ID>IN_2</ID>15 </input>
<input>
<ID>IN_3</ID>3 </input>
<output>
<ID>OUT</ID>254 </output>
<input>
<ID>SEL_0</ID>41 </input>
<input>
<ID>SEL_1</ID>258 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>533</ID>
<type>AA_LABEL</type>
<position>170.5,-129</position>
<gparam>LABEL_TEXT U2f</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>144</ID>
<type>AE_MUX_4x1</type>
<position>217,-127</position>
<input>
<ID>IN_0</ID>38 </input>
<input>
<ID>IN_1</ID>21 </input>
<input>
<ID>IN_2</ID>14 </input>
<input>
<ID>IN_3</ID>4 </input>
<output>
<ID>OUT</ID>253 </output>
<input>
<ID>SEL_0</ID>41 </input>
<input>
<ID>SEL_1</ID>258 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>534</ID>
<type>AA_LABEL</type>
<position>170.5,-133</position>
<gparam>LABEL_TEXT U2g</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>145</ID>
<type>AE_MUX_4x1</type>
<position>217,-141</position>
<input>
<ID>IN_0</ID>37 </input>
<input>
<ID>IN_1</ID>20 </input>
<input>
<ID>IN_2</ID>13 </input>
<input>
<ID>IN_3</ID>5 </input>
<output>
<ID>OUT</ID>252 </output>
<input>
<ID>SEL_0</ID>41 </input>
<input>
<ID>SEL_1</ID>258 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>535</ID>
<type>AA_LABEL</type>
<position>170.5,-137</position>
<gparam>LABEL_TEXT U2h</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>146</ID>
<type>AE_MUX_4x1</type>
<position>217,-155</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>19 </input>
<input>
<ID>IN_2</ID>12 </input>
<input>
<ID>IN_3</ID>6 </input>
<output>
<ID>OUT</ID>251 </output>
<input>
<ID>SEL_0</ID>41 </input>
<input>
<ID>SEL_1</ID>258 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>536</ID>
<type>AA_LABEL</type>
<position>170.5,-143</position>
<gparam>LABEL_TEXT U3a</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>147</ID>
<type>AE_MUX_4x1</type>
<position>217,-169</position>
<input>
<ID>IN_0</ID>35 </input>
<input>
<ID>IN_1</ID>18 </input>
<input>
<ID>IN_2</ID>11 </input>
<input>
<ID>IN_3</ID>7 </input>
<output>
<ID>OUT</ID>234 </output>
<input>
<ID>SEL_0</ID>41 </input>
<input>
<ID>SEL_1</ID>258 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>537</ID>
<type>AA_LABEL</type>
<position>170.5,-147</position>
<gparam>LABEL_TEXT U3b</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>538</ID>
<type>AA_LABEL</type>
<position>170.5,-151</position>
<gparam>LABEL_TEXT U3c</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>539</ID>
<type>AA_LABEL</type>
<position>170.5,-155</position>
<gparam>LABEL_TEXT U3d</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>540</ID>
<type>AA_LABEL</type>
<position>170.5,-159</position>
<gparam>LABEL_TEXT U3e</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>541</ID>
<type>AA_LABEL</type>
<position>170.5,-163</position>
<gparam>LABEL_TEXT U3f</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>542</ID>
<type>AA_LABEL</type>
<position>170.5,-167</position>
<gparam>LABEL_TEXT U3g</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>154</ID>
<type>AE_MUX_4x1</type>
<position>217,-183</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>17 </input>
<input>
<ID>IN_2</ID>10 </input>
<input>
<ID>IN_3</ID>8 </input>
<output>
<ID>OUT</ID>233 </output>
<input>
<ID>SEL_0</ID>41 </input>
<input>
<ID>SEL_1</ID>258 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>544</ID>
<type>AA_LABEL</type>
<position>170.5,-171</position>
<gparam>LABEL_TEXT U3h</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>546</ID>
<type>AA_LABEL</type>
<position>171,-177.5</position>
<gparam>LABEL_TEXT U4a</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>548</ID>
<type>AA_LABEL</type>
<position>171,-180.5</position>
<gparam>LABEL_TEXT U4b</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>550</ID>
<type>AA_LABEL</type>
<position>171,-183.5</position>
<gparam>LABEL_TEXT U4c</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>552</ID>
<type>AA_LABEL</type>
<position>171,-186.5</position>
<gparam>LABEL_TEXT U4d</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>163</ID>
<type>AE_SMALL_INVERTER</type>
<position>167.5,-239</position>
<input>
<ID>IN_0</ID>110 </input>
<output>
<ID>OUT_0</ID>170 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>164</ID>
<type>AE_SMALL_INVERTER</type>
<position>167.5,-231</position>
<input>
<ID>IN_0</ID>257 </input>
<output>
<ID>OUT_0</ID>169 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>554</ID>
<type>AA_LABEL</type>
<position>171,-189.5</position>
<gparam>LABEL_TEXT U4e</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>165</ID>
<type>AE_SMALL_INVERTER</type>
<position>167.5,-223</position>
<input>
<ID>IN_0</ID>63 </input>
<output>
<ID>OUT_0</ID>171 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>166</ID>
<type>AE_SMALL_INVERTER</type>
<position>167.5,-215</position>
<input>
<ID>IN_0</ID>61 </input>
<output>
<ID>OUT_0</ID>172 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>556</ID>
<type>AA_LABEL</type>
<position>171,-192.5</position>
<gparam>LABEL_TEXT U4f</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>558</ID>
<type>AA_LABEL</type>
<position>171,-195.5</position>
<gparam>LABEL_TEXT U4g</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>559</ID>
<type>AA_LABEL</type>
<position>171,-198.5</position>
<gparam>LABEL_TEXT U4h</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>584</ID>
<type>AA_LABEL</type>
<position>217,-77</position>
<gparam>LABEL_TEXT 74LS253</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>585</ID>
<type>AA_LABEL</type>
<position>217,-90</position>
<gparam>LABEL_TEXT U5a</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>586</ID>
<type>AA_LABEL</type>
<position>217,-104</position>
<gparam>LABEL_TEXT U5b</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>587</ID>
<type>AA_LABEL</type>
<position>217,-118</position>
<gparam>LABEL_TEXT U5c</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>588</ID>
<type>AA_LABEL</type>
<position>217,-132</position>
<gparam>LABEL_TEXT U5d</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>589</ID>
<type>AA_LABEL</type>
<position>217,-146</position>
<gparam>LABEL_TEXT U5e</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>590</ID>
<type>AA_LABEL</type>
<position>217,-160</position>
<gparam>LABEL_TEXT U5f</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>591</ID>
<type>AA_LABEL</type>
<position>217,-174</position>
<gparam>LABEL_TEXT U5g</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>592</ID>
<type>AA_LABEL</type>
<position>217,-188</position>
<gparam>LABEL_TEXT U5h</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>601</ID>
<type>AA_LABEL</type>
<position>151,-217</position>
<gparam>LABEL_TEXT U2i</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>602</ID>
<type>AA_LABEL</type>
<position>151,-225</position>
<gparam>LABEL_TEXT U2j</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>603</ID>
<type>AA_LABEL</type>
<position>151,-233</position>
<gparam>LABEL_TEXT U2k</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>604</ID>
<type>AA_LABEL</type>
<position>151,-241</position>
<gparam>LABEL_TEXT U2l</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>605</ID>
<type>AA_LABEL</type>
<position>151,-249</position>
<gparam>LABEL_TEXT U2m</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>606</ID>
<type>AA_LABEL</type>
<position>151,-257</position>
<gparam>LABEL_TEXT U2n</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>607</ID>
<type>AA_LABEL</type>
<position>151,-265</position>
<gparam>LABEL_TEXT U2o</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>608</ID>
<type>AA_LABEL</type>
<position>151,-273</position>
<gparam>LABEL_TEXT U2p</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>609</ID>
<type>AA_LABEL</type>
<position>164,-212</position>
<gparam>LABEL_TEXT U1i</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>610</ID>
<type>AA_LABEL</type>
<position>164,-216</position>
<gparam>LABEL_TEXT U1j</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>611</ID>
<type>AA_LABEL</type>
<position>164,-220</position>
<gparam>LABEL_TEXT U1k</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>612</ID>
<type>AA_LABEL</type>
<position>164,-224</position>
<gparam>LABEL_TEXT U1l</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>613</ID>
<type>AA_LABEL</type>
<position>164,-228</position>
<gparam>LABEL_TEXT U1m</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>614</ID>
<type>AA_LABEL</type>
<position>164,-232</position>
<gparam>LABEL_TEXT U1n</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>615</ID>
<type>AA_LABEL</type>
<position>164,-236</position>
<gparam>LABEL_TEXT U1o</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>616</ID>
<type>AA_LABEL</type>
<position>164,-240</position>
<gparam>LABEL_TEXT U1p</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>617</ID>
<type>AA_LABEL</type>
<position>164,-244</position>
<gparam>LABEL_TEXT U1q</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>618</ID>
<type>AA_LABEL</type>
<position>164,-248</position>
<gparam>LABEL_TEXT U1r</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>619</ID>
<type>AA_LABEL</type>
<position>164,-252</position>
<gparam>LABEL_TEXT U1s</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>620</ID>
<type>AA_LABEL</type>
<position>164,-256</position>
<gparam>LABEL_TEXT U1t</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>621</ID>
<type>AA_LABEL</type>
<position>164,-260</position>
<gparam>LABEL_TEXT U1u</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>622</ID>
<type>AA_LABEL</type>
<position>164,-264</position>
<gparam>LABEL_TEXT U1v</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>623</ID>
<type>AA_LABEL</type>
<position>164,-268</position>
<gparam>LABEL_TEXT U1w</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>624</ID>
<type>AA_LABEL</type>
<position>164,-272</position>
<gparam>LABEL_TEXT U1x</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>625</ID>
<type>AA_LABEL</type>
<position>132,-276</position>
<gparam>LABEL_TEXT 74HC283</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>626</ID>
<type>AA_LABEL</type>
<position>123,-276</position>
<gparam>LABEL_TEXT U6a</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>627</ID>
<type>AA_LABEL</type>
<position>141,-276</position>
<gparam>LABEL_TEXT U6b</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>628</ID>
<type>AA_LABEL</type>
<position>286,-105.5</position>
<gparam>LABEL_TEXT 74HC257</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>630</ID>
<type>AA_LABEL</type>
<position>286,-112.5</position>
<gparam>LABEL_TEXT U7a</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>631</ID>
<type>AA_LABEL</type>
<position>286,-119.5</position>
<gparam>LABEL_TEXT U7b</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>632</ID>
<type>AA_LABEL</type>
<position>286,-126.5</position>
<gparam>LABEL_TEXT U7c</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>633</ID>
<type>AA_LABEL</type>
<position>286,-133.5</position>
<gparam>LABEL_TEXT U7d</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>634</ID>
<type>AA_LABEL</type>
<position>286,-140</position>
<gparam>LABEL_TEXT U7e</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>635</ID>
<type>AA_LABEL</type>
<position>286,-147</position>
<gparam>LABEL_TEXT U7f</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>636</ID>
<type>AA_LABEL</type>
<position>286,-154</position>
<gparam>LABEL_TEXT U7g</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>637</ID>
<type>AA_LABEL</type>
<position>286,-161</position>
<gparam>LABEL_TEXT U7h</gparam>
<gparam>TEXT_HEIGHT 0.8</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>279</ID>
<type>AE_FULLADDER_4BIT</type>
<position>123,-281</position>
<input>
<ID>IN_0</ID>111 </input>
<input>
<ID>IN_1</ID>109 </input>
<input>
<ID>IN_2</ID>81 </input>
<input>
<ID>IN_3</ID>62 </input>
<input>
<ID>IN_B_0</ID>175 </input>
<input>
<ID>IN_B_1</ID>176 </input>
<input>
<ID>IN_B_2</ID>177 </input>
<input>
<ID>IN_B_3</ID>178 </input>
<output>
<ID>OUT_0</ID>264 </output>
<output>
<ID>OUT_1</ID>265 </output>
<output>
<ID>OUT_2</ID>266 </output>
<output>
<ID>OUT_3</ID>267 </output>
<input>
<ID>carry_in</ID>128 </input>
<output>
<ID>carry_out</ID>268 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>284</ID>
<type>AE_FULLADDER_4BIT</type>
<position>141,-281</position>
<input>
<ID>IN_0</ID>119 </input>
<input>
<ID>IN_1</ID>117 </input>
<input>
<ID>IN_2</ID>115 </input>
<input>
<ID>IN_3</ID>113 </input>
<input>
<ID>IN_B_0</ID>155 </input>
<input>
<ID>IN_B_1</ID>158 </input>
<input>
<ID>IN_B_2</ID>173 </input>
<input>
<ID>IN_B_3</ID>174 </input>
<output>
<ID>OUT_0</ID>260 </output>
<output>
<ID>OUT_1</ID>261 </output>
<output>
<ID>OUT_2</ID>262 </output>
<output>
<ID>OUT_3</ID>263 </output>
<input>
<ID>carry_in</ID>41 </input>
<output>
<ID>carry_out</ID>128 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>349</ID>
<type>AA_AND2</type>
<position>159.5,-244</position>
<input>
<ID>IN_0</ID>258 </input>
<input>
<ID>IN_1</ID>112 </input>
<output>
<ID>OUT</ID>146 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>350</ID>
<type>AA_AND2</type>
<position>159.5,-248</position>
<input>
<ID>IN_0</ID>259 </input>
<input>
<ID>IN_1</ID>163 </input>
<output>
<ID>OUT</ID>145 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>351</ID>
<type>AA_AND2</type>
<position>159.5,-252</position>
<input>
<ID>IN_0</ID>258 </input>
<input>
<ID>IN_1</ID>114 </input>
<output>
<ID>OUT</ID>144 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>352</ID>
<type>AA_AND2</type>
<position>159.5,-256</position>
<input>
<ID>IN_0</ID>259 </input>
<input>
<ID>IN_1</ID>161 </input>
<output>
<ID>OUT</ID>143 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>353</ID>
<type>AA_AND2</type>
<position>159.5,-260</position>
<input>
<ID>IN_0</ID>258 </input>
<input>
<ID>IN_1</ID>116 </input>
<output>
<ID>OUT</ID>142 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>354</ID>
<type>AA_AND2</type>
<position>159.5,-264</position>
<input>
<ID>IN_0</ID>259 </input>
<input>
<ID>IN_1</ID>159 </input>
<output>
<ID>OUT</ID>141 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>355</ID>
<type>AA_AND2</type>
<position>159.5,-268</position>
<input>
<ID>IN_0</ID>258 </input>
<input>
<ID>IN_1</ID>118 </input>
<output>
<ID>OUT</ID>139 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>356</ID>
<type>AA_AND2</type>
<position>159.5,-272</position>
<input>
<ID>IN_0</ID>259 </input>
<input>
<ID>IN_1</ID>157 </input>
<output>
<ID>OUT</ID>140 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>357</ID>
<type>AA_AND2</type>
<position>159.5,-212</position>
<input>
<ID>IN_0</ID>258 </input>
<input>
<ID>IN_1</ID>61 </input>
<output>
<ID>OUT</ID>154 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>358</ID>
<type>AA_AND2</type>
<position>159.5,-216</position>
<input>
<ID>IN_0</ID>259 </input>
<input>
<ID>IN_1</ID>172 </input>
<output>
<ID>OUT</ID>153 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>359</ID>
<type>AA_AND2</type>
<position>159.5,-220</position>
<input>
<ID>IN_0</ID>258 </input>
<input>
<ID>IN_1</ID>63 </input>
<output>
<ID>OUT</ID>152 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>360</ID>
<type>AA_AND2</type>
<position>159.5,-224</position>
<input>
<ID>IN_0</ID>259 </input>
<input>
<ID>IN_1</ID>171 </input>
<output>
<ID>OUT</ID>151 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>361</ID>
<type>AA_AND2</type>
<position>159.5,-228</position>
<input>
<ID>IN_0</ID>258 </input>
<input>
<ID>IN_1</ID>257 </input>
<output>
<ID>OUT</ID>150 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>362</ID>
<type>AA_AND2</type>
<position>159.5,-232</position>
<input>
<ID>IN_0</ID>259 </input>
<input>
<ID>IN_1</ID>169 </input>
<output>
<ID>OUT</ID>149 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>363</ID>
<type>AA_AND2</type>
<position>159.5,-236</position>
<input>
<ID>IN_0</ID>258 </input>
<input>
<ID>IN_1</ID>110 </input>
<output>
<ID>OUT</ID>148 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>364</ID>
<type>AA_AND2</type>
<position>159.5,-240</position>
<input>
<ID>IN_0</ID>259 </input>
<input>
<ID>IN_1</ID>170 </input>
<output>
<ID>OUT</ID>147 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>365</ID>
<type>AE_OR2</type>
<position>151,-270</position>
<input>
<ID>IN_0</ID>140 </input>
<input>
<ID>IN_1</ID>139 </input>
<output>
<ID>OUT</ID>155 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>366</ID>
<type>AE_OR2</type>
<position>151,-262</position>
<input>
<ID>IN_0</ID>141 </input>
<input>
<ID>IN_1</ID>142 </input>
<output>
<ID>OUT</ID>158 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>367</ID>
<type>AE_OR2</type>
<position>151,-254</position>
<input>
<ID>IN_0</ID>143 </input>
<input>
<ID>IN_1</ID>144 </input>
<output>
<ID>OUT</ID>173 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>368</ID>
<type>AE_OR2</type>
<position>151,-246</position>
<input>
<ID>IN_0</ID>145 </input>
<input>
<ID>IN_1</ID>146 </input>
<output>
<ID>OUT</ID>174 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>369</ID>
<type>AE_OR2</type>
<position>151,-238</position>
<input>
<ID>IN_0</ID>147 </input>
<input>
<ID>IN_1</ID>148 </input>
<output>
<ID>OUT</ID>175 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>370</ID>
<type>AE_OR2</type>
<position>151,-230</position>
<input>
<ID>IN_0</ID>149 </input>
<input>
<ID>IN_1</ID>150 </input>
<output>
<ID>OUT</ID>176 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>371</ID>
<type>AE_OR2</type>
<position>151,-222</position>
<input>
<ID>IN_0</ID>151 </input>
<input>
<ID>IN_1</ID>152 </input>
<output>
<ID>OUT</ID>177 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>372</ID>
<type>AE_OR2</type>
<position>151,-214</position>
<input>
<ID>IN_0</ID>153 </input>
<input>
<ID>IN_1</ID>154 </input>
<output>
<ID>OUT</ID>178 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>373</ID>
<type>AE_SMALL_INVERTER</type>
<position>167.5,-271</position>
<input>
<ID>IN_0</ID>118 </input>
<output>
<ID>OUT_0</ID>157 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>374</ID>
<type>AE_SMALL_INVERTER</type>
<position>167.5,-263</position>
<input>
<ID>IN_0</ID>116 </input>
<output>
<ID>OUT_0</ID>159 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>375</ID>
<type>AE_SMALL_INVERTER</type>
<position>167.5,-255</position>
<input>
<ID>IN_0</ID>114 </input>
<output>
<ID>OUT_0</ID>161 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>376</ID>
<type>AE_SMALL_INVERTER</type>
<position>167.5,-247</position>
<input>
<ID>IN_0</ID>112 </input>
<output>
<ID>OUT_0</ID>163 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>378</ID>
<type>AA_MUX_2x1</type>
<position>286,-131</position>
<input>
<ID>IN_0</ID>264 </input>
<input>
<ID>IN_1</ID>253 </input>
<output>
<ID>OUT</ID>184 </output>
<input>
<ID>SEL_0</ID>256 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>379</ID>
<type>AA_MUX_2x1</type>
<position>286,-124</position>
<input>
<ID>IN_0</ID>265 </input>
<input>
<ID>IN_1</ID>254 </input>
<output>
<ID>OUT</ID>183 </output>
<input>
<ID>SEL_0</ID>256 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>380</ID>
<type>AA_MUX_2x1</type>
<position>286,-117</position>
<input>
<ID>IN_0</ID>266 </input>
<input>
<ID>IN_1</ID>255 </input>
<output>
<ID>OUT</ID>182 </output>
<input>
<ID>SEL_0</ID>256 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>381</ID>
<type>AA_MUX_2x1</type>
<position>286,-110</position>
<input>
<ID>IN_0</ID>267 </input>
<input>
<ID>IN_1</ID>219 </input>
<output>
<ID>OUT</ID>181 </output>
<input>
<ID>SEL_0</ID>256 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>382</ID>
<type>AA_MUX_2x1</type>
<position>286,-158.5</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>233 </input>
<output>
<ID>OUT</ID>188 </output>
<input>
<ID>SEL_0</ID>256 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>383</ID>
<type>AA_MUX_2x1</type>
<position>286,-151.5</position>
<input>
<ID>IN_0</ID>261 </input>
<input>
<ID>IN_1</ID>234 </input>
<output>
<ID>OUT</ID>187 </output>
<input>
<ID>SEL_0</ID>256 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>384</ID>
<type>AA_MUX_2x1</type>
<position>286,-144.5</position>
<input>
<ID>IN_0</ID>262 </input>
<input>
<ID>IN_1</ID>251 </input>
<output>
<ID>OUT</ID>186 </output>
<input>
<ID>SEL_0</ID>256 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>385</ID>
<type>AA_MUX_2x1</type>
<position>286,-137.5</position>
<input>
<ID>IN_0</ID>263 </input>
<input>
<ID>IN_1</ID>252 </input>
<output>
<ID>OUT</ID>185 </output>
<input>
<ID>SEL_0</ID>256 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>386</ID>
<type>AA_LABEL</type>
<position>302,-136</position>
<gparam>LABEL_TEXT G3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>387</ID>
<type>AA_LABEL</type>
<position>302,-140</position>
<gparam>LABEL_TEXT G2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>388</ID>
<type>AA_LABEL</type>
<position>302,-144</position>
<gparam>LABEL_TEXT G1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>205,-177,205,-82</points>
<intersection>-177 2</intersection>
<intersection>-82 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>205,-82,214,-82</points>
<connection>
<GID>141</GID>
<name>IN_3</name></connection>
<intersection>205 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>177,-177,205,-177</points>
<connection>
<GID>131</GID>
<name>OUT_0</name></connection>
<intersection>205 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>206,-180,206,-96</points>
<intersection>-180 2</intersection>
<intersection>-96 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>206,-96,214,-96</points>
<connection>
<GID>142</GID>
<name>IN_3</name></connection>
<intersection>206 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>177,-180,206,-180</points>
<connection>
<GID>132</GID>
<name>OUT_0</name></connection>
<intersection>206 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207,-183,207,-110</points>
<intersection>-183 2</intersection>
<intersection>-110 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>207,-110,214,-110</points>
<connection>
<GID>143</GID>
<name>IN_3</name></connection>
<intersection>207 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>177,-183,207,-183</points>
<connection>
<GID>133</GID>
<name>OUT_0</name></connection>
<intersection>207 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>208,-186,208,-124</points>
<intersection>-186 2</intersection>
<intersection>-124 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>208,-124,214,-124</points>
<connection>
<GID>144</GID>
<name>IN_3</name></connection>
<intersection>208 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>177,-186,208,-186</points>
<connection>
<GID>134</GID>
<name>OUT_0</name></connection>
<intersection>208 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>209,-189,209,-138</points>
<intersection>-189 2</intersection>
<intersection>-138 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>209,-138,214,-138</points>
<connection>
<GID>145</GID>
<name>IN_3</name></connection>
<intersection>209 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>177,-189,209,-189</points>
<connection>
<GID>135</GID>
<name>OUT_0</name></connection>
<intersection>209 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>210,-192,210,-152</points>
<intersection>-192 2</intersection>
<intersection>-152 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>210,-152,214,-152</points>
<connection>
<GID>146</GID>
<name>IN_3</name></connection>
<intersection>210 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>177,-192,210,-192</points>
<connection>
<GID>136</GID>
<name>OUT_0</name></connection>
<intersection>210 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>211,-195,211,-166</points>
<intersection>-195 2</intersection>
<intersection>-166 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>211,-166,214,-166</points>
<connection>
<GID>147</GID>
<name>IN_3</name></connection>
<intersection>211 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>177,-195,211,-195</points>
<connection>
<GID>137</GID>
<name>OUT_0</name></connection>
<intersection>211 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>212,-198,212,-180</points>
<intersection>-198 2</intersection>
<intersection>-180 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>212,-180,214,-180</points>
<connection>
<GID>154</GID>
<name>IN_3</name></connection>
<intersection>212 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>177,-198,212,-198</points>
<connection>
<GID>140</GID>
<name>OUT_0</name></connection>
<intersection>212 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>196,-143,196,-84</points>
<intersection>-143 2</intersection>
<intersection>-84 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>196,-84,214,-84</points>
<connection>
<GID>141</GID>
<name>IN_2</name></connection>
<intersection>196 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>178.5,-143,196,-143</points>
<connection>
<GID>123</GID>
<name>OUT</name></connection>
<intersection>196 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-182,201,-171</points>
<intersection>-182 1</intersection>
<intersection>-171 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>201,-182,214,-182</points>
<connection>
<GID>154</GID>
<name>IN_2</name></connection>
<intersection>201 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>178.5,-171,201,-171</points>
<connection>
<GID>130</GID>
<name>OUT</name></connection>
<intersection>201 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-168,201,-167</points>
<intersection>-168 1</intersection>
<intersection>-167 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>201,-168,214,-168</points>
<connection>
<GID>147</GID>
<name>IN_2</name></connection>
<intersection>201 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>178.5,-167,201,-167</points>
<connection>
<GID>129</GID>
<name>OUT</name></connection>
<intersection>201 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>201,-163,201,-154</points>
<intersection>-163 2</intersection>
<intersection>-154 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>201,-154,214,-154</points>
<connection>
<GID>146</GID>
<name>IN_2</name></connection>
<intersection>201 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>178.5,-163,201,-163</points>
<connection>
<GID>128</GID>
<name>OUT</name></connection>
<intersection>201 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>200,-159,200,-140</points>
<intersection>-159 2</intersection>
<intersection>-140 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>200,-140,214,-140</points>
<connection>
<GID>145</GID>
<name>IN_2</name></connection>
<intersection>200 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>178.5,-159,200,-159</points>
<connection>
<GID>127</GID>
<name>OUT</name></connection>
<intersection>200 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>199,-155,199,-126</points>
<intersection>-155 2</intersection>
<intersection>-126 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>199,-126,214,-126</points>
<connection>
<GID>144</GID>
<name>IN_2</name></connection>
<intersection>199 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>178.5,-155,199,-155</points>
<connection>
<GID>126</GID>
<name>OUT</name></connection>
<intersection>199 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>198,-151,198,-112</points>
<intersection>-151 2</intersection>
<intersection>-112 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>198,-112,214,-112</points>
<connection>
<GID>143</GID>
<name>IN_2</name></connection>
<intersection>198 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>178.5,-151,198,-151</points>
<connection>
<GID>125</GID>
<name>OUT</name></connection>
<intersection>198 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>197,-147,197,-98</points>
<intersection>-147 2</intersection>
<intersection>-98 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>197,-98,214,-98</points>
<connection>
<GID>142</GID>
<name>IN_2</name></connection>
<intersection>197 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>178.5,-147,197,-147</points>
<connection>
<GID>124</GID>
<name>OUT</name></connection>
<intersection>197 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>188,-184,188,-137</points>
<intersection>-184 1</intersection>
<intersection>-137 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>188,-184,214,-184</points>
<connection>
<GID>154</GID>
<name>IN_1</name></connection>
<intersection>188 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>178,-137,188,-137</points>
<connection>
<GID>122</GID>
<name>OUT</name></connection>
<intersection>188 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189,-170,189,-133</points>
<intersection>-170 1</intersection>
<intersection>-133 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189,-170,214,-170</points>
<connection>
<GID>147</GID>
<name>IN_1</name></connection>
<intersection>189 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>178,-133,189,-133</points>
<connection>
<GID>121</GID>
<name>OUT</name></connection>
<intersection>189 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>190,-156,190,-129</points>
<intersection>-156 1</intersection>
<intersection>-129 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>190,-156,214,-156</points>
<connection>
<GID>146</GID>
<name>IN_1</name></connection>
<intersection>190 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>178,-129,190,-129</points>
<connection>
<GID>120</GID>
<name>OUT</name></connection>
<intersection>190 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191,-142,191,-125</points>
<intersection>-142 1</intersection>
<intersection>-125 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191,-142,214,-142</points>
<connection>
<GID>145</GID>
<name>IN_1</name></connection>
<intersection>191 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>178,-125,191,-125</points>
<connection>
<GID>119</GID>
<name>OUT</name></connection>
<intersection>191 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>192,-128,192,-121</points>
<intersection>-128 1</intersection>
<intersection>-121 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>192,-128,214,-128</points>
<connection>
<GID>144</GID>
<name>IN_1</name></connection>
<intersection>192 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>178,-121,192,-121</points>
<connection>
<GID>118</GID>
<name>OUT</name></connection>
<intersection>192 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>192,-117,192,-114</points>
<intersection>-117 2</intersection>
<intersection>-114 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>192,-114,214,-114</points>
<connection>
<GID>143</GID>
<name>IN_1</name></connection>
<intersection>192 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>178,-117,192,-117</points>
<connection>
<GID>117</GID>
<name>OUT</name></connection>
<intersection>192 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>192,-113,192,-100</points>
<intersection>-113 2</intersection>
<intersection>-100 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>192,-100,214,-100</points>
<connection>
<GID>142</GID>
<name>IN_1</name></connection>
<intersection>192 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>178,-113,192,-113</points>
<connection>
<GID>116</GID>
<name>OUT</name></connection>
<intersection>192 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191,-109,191,-86</points>
<intersection>-109 2</intersection>
<intersection>-86 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191,-86,214,-86</points>
<connection>
<GID>141</GID>
<name>IN_1</name></connection>
<intersection>191 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>178,-109,191,-109</points>
<connection>
<GID>115</GID>
<name>OUT</name></connection>
<intersection>191 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187,-88,187,-75</points>
<intersection>-88 1</intersection>
<intersection>-75 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>187,-88,214,-88</points>
<connection>
<GID>141</GID>
<name>IN_0</name></connection>
<intersection>187 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>178,-75,187,-75</points>
<connection>
<GID>89</GID>
<name>OUT</name></connection>
<intersection>187 0</intersection></hsegment></shape></wire>
<wire>
<ID>219</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>259,-109,259,-85</points>
<intersection>-109 1</intersection>
<intersection>-85 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>259,-109,284,-109</points>
<connection>
<GID>381</GID>
<name>IN_1</name></connection>
<intersection>259 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220,-85,259,-85</points>
<connection>
<GID>141</GID>
<name>OUT</name></connection>
<intersection>259 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>180,-186,180,-103</points>
<intersection>-186 1</intersection>
<intersection>-103 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>180,-186,214,-186</points>
<connection>
<GID>154</GID>
<name>IN_0</name></connection>
<intersection>180 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>178,-103,180,-103</points>
<connection>
<GID>114</GID>
<name>OUT</name></connection>
<intersection>180 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>181,-172,181,-99</points>
<intersection>-172 1</intersection>
<intersection>-99 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>181,-172,214,-172</points>
<connection>
<GID>147</GID>
<name>IN_0</name></connection>
<intersection>181 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>178,-99,181,-99</points>
<connection>
<GID>113</GID>
<name>OUT</name></connection>
<intersection>181 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>182,-158,182,-95</points>
<intersection>-158 1</intersection>
<intersection>-95 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>182,-158,214,-158</points>
<connection>
<GID>146</GID>
<name>IN_0</name></connection>
<intersection>182 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>178,-95,182,-95</points>
<connection>
<GID>112</GID>
<name>OUT</name></connection>
<intersection>182 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>183,-144,183,-91</points>
<intersection>-144 1</intersection>
<intersection>-91 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>183,-144,214,-144</points>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<intersection>183 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>178,-91,183,-91</points>
<connection>
<GID>111</GID>
<name>OUT</name></connection>
<intersection>183 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184,-130,184,-87</points>
<intersection>-130 1</intersection>
<intersection>-87 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>184,-130,214,-130</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>178,-87,184,-87</points>
<connection>
<GID>110</GID>
<name>OUT</name></connection>
<intersection>184 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185,-116,185,-83</points>
<intersection>-116 1</intersection>
<intersection>-83 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>185,-116,214,-116</points>
<connection>
<GID>143</GID>
<name>IN_0</name></connection>
<intersection>185 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>178,-83,185,-83</points>
<connection>
<GID>109</GID>
<name>OUT</name></connection>
<intersection>185 0</intersection></hsegment></shape></wire>
<wire>
<ID>233</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>259,-183,259,-157.5</points>
<intersection>-183 2</intersection>
<intersection>-157.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>259,-157.5,284,-157.5</points>
<connection>
<GID>382</GID>
<name>IN_1</name></connection>
<intersection>259 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220,-183,259,-183</points>
<connection>
<GID>154</GID>
<name>OUT</name></connection>
<intersection>259 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>186,-102,186,-79</points>
<intersection>-102 1</intersection>
<intersection>-79 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>186,-102,214,-102</points>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<intersection>186 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>178,-79,186,-79</points>
<connection>
<GID>91</GID>
<name>OUT</name></connection>
<intersection>186 0</intersection></hsegment></shape></wire>
<wire>
<ID>234</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>257,-169,257,-150.5</points>
<intersection>-169 2</intersection>
<intersection>-150.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>257,-150.5,284,-150.5</points>
<connection>
<GID>383</GID>
<name>IN_1</name></connection>
<intersection>257 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220,-169,257,-169</points>
<connection>
<GID>147</GID>
<name>OUT</name></connection>
<intersection>257 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>234.5,-280,234.5,-68</points>
<connection>
<GID>81</GID>
<name>OUT_0</name></connection>
<intersection>-280 22</intersection>
<intersection>-178 3</intersection>
<intersection>-164 4</intersection>
<intersection>-150 7</intersection>
<intersection>-136 8</intersection>
<intersection>-122 9</intersection>
<intersection>-108 10</intersection>
<intersection>-94 11</intersection>
<intersection>-80 12</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>218,-178,234.5,-178</points>
<connection>
<GID>154</GID>
<name>SEL_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>218,-164,234.5,-164</points>
<connection>
<GID>147</GID>
<name>SEL_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>218,-150,234.5,-150</points>
<connection>
<GID>146</GID>
<name>SEL_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>218,-136,234.5,-136</points>
<connection>
<GID>145</GID>
<name>SEL_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>218,-122,234.5,-122</points>
<connection>
<GID>144</GID>
<name>SEL_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>218,-108,234.5,-108</points>
<connection>
<GID>143</GID>
<name>SEL_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>218,-94,234.5,-94</points>
<connection>
<GID>142</GID>
<name>SEL_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>218,-80,234.5,-80</points>
<connection>
<GID>141</GID>
<name>SEL_0</name></connection>
<intersection>234.5 0</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>149,-280,234.5,-280</points>
<connection>
<GID>284</GID>
<name>carry_in</name></connection>
<intersection>234.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>251</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>255,-155,255,-143.5</points>
<intersection>-155 2</intersection>
<intersection>-143.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>255,-143.5,284,-143.5</points>
<connection>
<GID>384</GID>
<name>IN_1</name></connection>
<intersection>255 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220,-155,255,-155</points>
<connection>
<GID>146</GID>
<name>OUT</name></connection>
<intersection>255 0</intersection></hsegment></shape></wire>
<wire>
<ID>252</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>253,-141,253,-136.5</points>
<intersection>-141 2</intersection>
<intersection>-136.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>253,-136.5,284,-136.5</points>
<connection>
<GID>385</GID>
<name>IN_1</name></connection>
<intersection>253 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220,-141,253,-141</points>
<connection>
<GID>145</GID>
<name>OUT</name></connection>
<intersection>253 0</intersection></hsegment></shape></wire>
<wire>
<ID>253</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>253,-130,253,-127</points>
<intersection>-130 3</intersection>
<intersection>-127 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>220,-127,253,-127</points>
<connection>
<GID>144</GID>
<name>OUT</name></connection>
<intersection>253 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>253,-130,284,-130</points>
<connection>
<GID>378</GID>
<name>IN_1</name></connection>
<intersection>253 0</intersection></hsegment></shape></wire>
<wire>
<ID>254</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>255,-123,255,-113</points>
<intersection>-123 1</intersection>
<intersection>-113 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>255,-123,284,-123</points>
<connection>
<GID>379</GID>
<name>IN_1</name></connection>
<intersection>255 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220,-113,255,-113</points>
<connection>
<GID>143</GID>
<name>OUT</name></connection>
<intersection>255 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148,-208,148,-68</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<intersection>-208 5</intersection>
<intersection>-142 1</intersection>
<intersection>-108 2</intersection>
<intersection>-74 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>148,-142,172.5,-142</points>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<intersection>148 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>148,-108,172,-108</points>
<connection>
<GID>115</GID>
<name>IN_0</name></connection>
<intersection>148 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>148,-74,172,-74</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<intersection>148 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>148,-208,169.5,-208</points>
<intersection>148 0</intersection>
<intersection>169.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>169.5,-215,169.5,-208</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<intersection>-211 7</intersection>
<intersection>-208 5</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>162.5,-211,169.5,-211</points>
<connection>
<GID>357</GID>
<name>IN_1</name></connection>
<intersection>169.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>255</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>257,-116,257,-99</points>
<intersection>-116 1</intersection>
<intersection>-99 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>257,-116,284,-116</points>
<connection>
<GID>380</GID>
<name>IN_1</name></connection>
<intersection>257 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>220,-99,257,-99</points>
<connection>
<GID>142</GID>
<name>OUT</name></connection>
<intersection>257 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118,-277,118,-68</points>
<connection>
<GID>71</GID>
<name>OUT_0</name></connection>
<connection>
<GID>279</GID>
<name>IN_3</name></connection>
<intersection>-177 7</intersection>
<intersection>-144 1</intersection>
<intersection>-110 3</intersection>
<intersection>-76 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>118,-144,172.5,-144</points>
<connection>
<GID>123</GID>
<name>IN_1</name></connection>
<intersection>118 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>118,-110,172,-110</points>
<connection>
<GID>115</GID>
<name>IN_1</name></connection>
<intersection>118 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>118,-76,172,-76</points>
<connection>
<GID>89</GID>
<name>IN_1</name></connection>
<intersection>118 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>118,-177,173,-177</points>
<connection>
<GID>131</GID>
<name>IN_0</name></connection>
<intersection>118 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-207,151,-68</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>-207 5</intersection>
<intersection>-146 1</intersection>
<intersection>-112 2</intersection>
<intersection>-78 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>151,-146,172.5,-146</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>151,-112,172,-112</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>151,-78,172,-78</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>151,-207,172.5,-207</points>
<intersection>151 0</intersection>
<intersection>172.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>172.5,-223,172.5,-207</points>
<intersection>-223 7</intersection>
<intersection>-207 5</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>169.5,-223,172.5,-223</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<intersection>169.5 8</intersection>
<intersection>172.5 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>169.5,-223,169.5,-219</points>
<intersection>-223 7</intersection>
<intersection>-219 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>162.5,-219,169.5,-219</points>
<connection>
<GID>359</GID>
<name>IN_1</name></connection>
<intersection>169.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>256</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>290,-156,290,-73</points>
<intersection>-156 3</intersection>
<intersection>-149 4</intersection>
<intersection>-142 5</intersection>
<intersection>-135 6</intersection>
<intersection>-128.5 7</intersection>
<intersection>-121.5 8</intersection>
<intersection>-114.5 9</intersection>
<intersection>-107.5 10</intersection>
<intersection>-73 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>225.5,-73,225.5,-68</points>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection>
<intersection>-73 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>225.5,-73,290,-73</points>
<intersection>225.5 1</intersection>
<intersection>290 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>286,-156,290,-156</points>
<connection>
<GID>382</GID>
<name>SEL_0</name></connection>
<intersection>290 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>286,-149,290,-149</points>
<connection>
<GID>383</GID>
<name>SEL_0</name></connection>
<intersection>290 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>286,-142,290,-142</points>
<connection>
<GID>384</GID>
<name>SEL_0</name></connection>
<intersection>290 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>286,-135,290,-135</points>
<connection>
<GID>385</GID>
<name>SEL_0</name></connection>
<intersection>290 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>286,-128.5,290,-128.5</points>
<connection>
<GID>378</GID>
<name>SEL_0</name></connection>
<intersection>290 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>286,-121.5,290,-121.5</points>
<connection>
<GID>379</GID>
<name>SEL_0</name></connection>
<intersection>290 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>286,-114.5,290,-114.5</points>
<connection>
<GID>380</GID>
<name>SEL_0</name></connection>
<intersection>290 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>286,-107.5,290,-107.5</points>
<connection>
<GID>381</GID>
<name>SEL_0</name></connection>
<intersection>290 0</intersection></hsegment></shape></wire>
<wire>
<ID>257</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>154,-206,154,-68</points>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection>
<intersection>-206 1</intersection>
<intersection>-150 8</intersection>
<intersection>-116 6</intersection>
<intersection>-82 7</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>154,-206,175.5,-206</points>
<intersection>154 0</intersection>
<intersection>175.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>175.5,-231,175.5,-206</points>
<intersection>-231 3</intersection>
<intersection>-206 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>169.5,-231,175.5,-231</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<intersection>169.5 4</intersection>
<intersection>175.5 2</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>169.5,-231,169.5,-227</points>
<intersection>-231 3</intersection>
<intersection>-227 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>162.5,-227,169.5,-227</points>
<connection>
<GID>361</GID>
<name>IN_1</name></connection>
<intersection>169.5 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>154,-116,172,-116</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<intersection>154 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>154,-82,172,-82</points>
<connection>
<GID>109</GID>
<name>IN_0</name></connection>
<intersection>154 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>154,-150,172.5,-150</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<intersection>154 0</intersection></hsegment></shape></wire>
<wire>
<ID>258</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>196.5,-269,196.5,-213</points>
<intersection>-269 1</intersection>
<intersection>-261 5</intersection>
<intersection>-253 7</intersection>
<intersection>-245 9</intersection>
<intersection>-241 2</intersection>
<intersection>-237 17</intersection>
<intersection>-229 15</intersection>
<intersection>-221 13</intersection>
<intersection>-213 11</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>162.5,-269,196.5,-269</points>
<connection>
<GID>355</GID>
<name>IN_0</name></connection>
<intersection>196.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>196.5,-241,231.5,-241</points>
<intersection>196.5 0</intersection>
<intersection>231.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>231.5,-241,231.5,-68</points>
<connection>
<GID>80</GID>
<name>OUT_0</name></connection>
<intersection>-241 2</intersection>
<intersection>-177 22</intersection>
<intersection>-163 26</intersection>
<intersection>-149 31</intersection>
<intersection>-135 36</intersection>
<intersection>-121 41</intersection>
<intersection>-107 46</intersection>
<intersection>-93 51</intersection>
<intersection>-79 52</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>162.5,-261,196.5,-261</points>
<connection>
<GID>353</GID>
<name>IN_0</name></connection>
<intersection>196.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>162.5,-253,196.5,-253</points>
<connection>
<GID>351</GID>
<name>IN_0</name></connection>
<intersection>196.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>162.5,-245,196.5,-245</points>
<connection>
<GID>349</GID>
<name>IN_0</name></connection>
<intersection>196.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>162.5,-213,196.5,-213</points>
<connection>
<GID>357</GID>
<name>IN_0</name></connection>
<intersection>196.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>162.5,-221,196.5,-221</points>
<connection>
<GID>359</GID>
<name>IN_0</name></connection>
<intersection>196.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>162.5,-229,196.5,-229</points>
<connection>
<GID>361</GID>
<name>IN_0</name></connection>
<intersection>196.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>162.5,-237,196.5,-237</points>
<connection>
<GID>363</GID>
<name>IN_0</name></connection>
<intersection>196.5 0</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>217,-177,231.5,-177</points>
<intersection>217 24</intersection>
<intersection>231.5 3</intersection></hsegment>
<vsegment>
<ID>24</ID>
<points>217,-178,217,-177</points>
<connection>
<GID>154</GID>
<name>SEL_1</name></connection>
<intersection>-177 22</intersection></vsegment>
<hsegment>
<ID>26</ID>
<points>217,-163,231.5,-163</points>
<intersection>217 29</intersection>
<intersection>231.5 3</intersection></hsegment>
<vsegment>
<ID>29</ID>
<points>217,-164,217,-163</points>
<connection>
<GID>147</GID>
<name>SEL_1</name></connection>
<intersection>-163 26</intersection></vsegment>
<hsegment>
<ID>31</ID>
<points>217,-149,231.5,-149</points>
<intersection>217 33</intersection>
<intersection>231.5 3</intersection></hsegment>
<vsegment>
<ID>33</ID>
<points>217,-150,217,-149</points>
<connection>
<GID>146</GID>
<name>SEL_1</name></connection>
<intersection>-149 31</intersection></vsegment>
<hsegment>
<ID>36</ID>
<points>217,-135,231.5,-135</points>
<intersection>217 38</intersection>
<intersection>231.5 3</intersection></hsegment>
<vsegment>
<ID>38</ID>
<points>217,-136,217,-135</points>
<connection>
<GID>145</GID>
<name>SEL_1</name></connection>
<intersection>-135 36</intersection></vsegment>
<hsegment>
<ID>41</ID>
<points>217,-121,231.5,-121</points>
<intersection>217 43</intersection>
<intersection>231.5 3</intersection></hsegment>
<vsegment>
<ID>43</ID>
<points>217,-122,217,-121</points>
<connection>
<GID>144</GID>
<name>SEL_1</name></connection>
<intersection>-121 41</intersection></vsegment>
<hsegment>
<ID>46</ID>
<points>217,-107,231.5,-107</points>
<intersection>217 48</intersection>
<intersection>231.5 3</intersection></hsegment>
<vsegment>
<ID>48</ID>
<points>217,-108,217,-107</points>
<connection>
<GID>143</GID>
<name>SEL_1</name></connection>
<intersection>-107 46</intersection></vsegment>
<hsegment>
<ID>51</ID>
<points>217,-93,231.5,-93</points>
<intersection>217 54</intersection>
<intersection>231.5 3</intersection></hsegment>
<hsegment>
<ID>52</ID>
<points>217,-79,231.5,-79</points>
<intersection>217 53</intersection>
<intersection>231.5 3</intersection></hsegment>
<vsegment>
<ID>53</ID>
<points>217,-80,217,-79</points>
<connection>
<GID>141</GID>
<name>SEL_1</name></connection>
<intersection>-79 52</intersection></vsegment>
<vsegment>
<ID>54</ID>
<points>217,-94,217,-93</points>
<connection>
<GID>142</GID>
<name>SEL_1</name></connection>
<intersection>-93 51</intersection></vsegment></shape></wire>
<wire>
<ID>259</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>193.5,-273,193.5,-217</points>
<intersection>-273 1</intersection>
<intersection>-265 16</intersection>
<intersection>-257 14</intersection>
<intersection>-249 12</intersection>
<intersection>-244 2</intersection>
<intersection>-241 10</intersection>
<intersection>-233 8</intersection>
<intersection>-225 6</intersection>
<intersection>-217 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>162.5,-273,193.5,-273</points>
<connection>
<GID>356</GID>
<name>IN_0</name></connection>
<intersection>193.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>193.5,-244,228.5,-244</points>
<intersection>193.5 0</intersection>
<intersection>228.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>228.5,-244,228.5,-68</points>
<connection>
<GID>79</GID>
<name>OUT_0</name></connection>
<intersection>-244 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>162.5,-217,193.5,-217</points>
<connection>
<GID>358</GID>
<name>IN_0</name></connection>
<intersection>193.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>162.5,-225,193.5,-225</points>
<connection>
<GID>360</GID>
<name>IN_0</name></connection>
<intersection>193.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>162.5,-233,193.5,-233</points>
<connection>
<GID>362</GID>
<name>IN_0</name></connection>
<intersection>193.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>162.5,-241,193.5,-241</points>
<connection>
<GID>364</GID>
<name>IN_0</name></connection>
<intersection>193.5 0</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>162.5,-249,193.5,-249</points>
<connection>
<GID>350</GID>
<name>IN_0</name></connection>
<intersection>193.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>162.5,-257,193.5,-257</points>
<connection>
<GID>352</GID>
<name>IN_0</name></connection>
<intersection>193.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>162.5,-265,193.5,-265</points>
<connection>
<GID>354</GID>
<name>IN_0</name></connection>
<intersection>193.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>260</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>282,-285,282,-159.5</points>
<intersection>-285 2</intersection>
<intersection>-159.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>282,-159.5,284,-159.5</points>
<connection>
<GID>382</GID>
<name>IN_0</name></connection>
<intersection>282 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>142.5,-285,282,-285</points>
<connection>
<GID>284</GID>
<name>OUT_0</name></connection>
<intersection>282 0</intersection></hsegment></shape></wire>
<wire>
<ID>261</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>281,-286,281,-152.5</points>
<intersection>-286 2</intersection>
<intersection>-152.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>281,-152.5,284,-152.5</points>
<connection>
<GID>383</GID>
<name>IN_0</name></connection>
<intersection>281 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>141.5,-286,281,-286</points>
<intersection>141.5 3</intersection>
<intersection>281 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>141.5,-286,141.5,-285</points>
<connection>
<GID>284</GID>
<name>OUT_1</name></connection>
<intersection>-286 2</intersection></vsegment></shape></wire>
<wire>
<ID>262</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>280,-287,280,-145.5</points>
<intersection>-287 2</intersection>
<intersection>-145.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>280,-145.5,284,-145.5</points>
<connection>
<GID>384</GID>
<name>IN_0</name></connection>
<intersection>280 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>140.5,-287,280,-287</points>
<intersection>140.5 3</intersection>
<intersection>280 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>140.5,-287,140.5,-285</points>
<connection>
<GID>284</GID>
<name>OUT_2</name></connection>
<intersection>-287 2</intersection></vsegment></shape></wire>
<wire>
<ID>263</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>279,-288,279,-138.5</points>
<intersection>-288 2</intersection>
<intersection>-138.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>279,-138.5,284,-138.5</points>
<connection>
<GID>385</GID>
<name>IN_0</name></connection>
<intersection>279 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>139.5,-288,279,-288</points>
<intersection>139.5 3</intersection>
<intersection>279 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>139.5,-288,139.5,-285</points>
<connection>
<GID>284</GID>
<name>OUT_3</name></connection>
<intersection>-288 2</intersection></vsegment></shape></wire>
<wire>
<ID>264</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>278,-289,278,-132</points>
<intersection>-289 2</intersection>
<intersection>-132 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>278,-132,284,-132</points>
<connection>
<GID>378</GID>
<name>IN_0</name></connection>
<intersection>278 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>124.5,-289,278,-289</points>
<intersection>124.5 3</intersection>
<intersection>278 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>124.5,-289,124.5,-285</points>
<connection>
<GID>279</GID>
<name>OUT_0</name></connection>
<intersection>-289 2</intersection></vsegment></shape></wire>
<wire>
<ID>265</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>277,-290,277,-125</points>
<intersection>-290 2</intersection>
<intersection>-125 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>277,-125,284,-125</points>
<connection>
<GID>379</GID>
<name>IN_0</name></connection>
<intersection>277 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>123.5,-290,277,-290</points>
<intersection>123.5 3</intersection>
<intersection>277 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>123.5,-290,123.5,-285</points>
<connection>
<GID>279</GID>
<name>OUT_1</name></connection>
<intersection>-290 2</intersection></vsegment></shape></wire>
<wire>
<ID>266</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>276,-291,276,-118</points>
<intersection>-291 2</intersection>
<intersection>-118 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>276,-118,284,-118</points>
<connection>
<GID>380</GID>
<name>IN_0</name></connection>
<intersection>276 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>122.5,-291,276,-291</points>
<intersection>122.5 3</intersection>
<intersection>276 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>122.5,-291,122.5,-285</points>
<connection>
<GID>279</GID>
<name>OUT_2</name></connection>
<intersection>-291 2</intersection></vsegment></shape></wire>
<wire>
<ID>267</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>275,-292,275,-111</points>
<intersection>-292 2</intersection>
<intersection>-111 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>275,-111,284,-111</points>
<connection>
<GID>381</GID>
<name>IN_0</name></connection>
<intersection>275 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>121.5,-292,275,-292</points>
<intersection>121.5 3</intersection>
<intersection>275 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>121.5,-292,121.5,-285</points>
<connection>
<GID>279</GID>
<name>OUT_3</name></connection>
<intersection>-292 2</intersection></vsegment></shape></wire>
<wire>
<ID>268</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>114,-293,305,-293</points>
<intersection>114 4</intersection>
<intersection>305 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>305,-293,305,-114</points>
<intersection>-293 1</intersection>
<intersection>-114 6</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>114,-293,114,-280</points>
<intersection>-293 1</intersection>
<intersection>-280 7</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>300.5,-114,305,-114</points>
<connection>
<GID>404</GID>
<name>N_in1</name></connection>
<intersection>305 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>114,-280,115,-280</points>
<connection>
<GID>279</GID>
<name>carry_out</name></connection>
<intersection>114 4</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121,-204,121,-68</points>
<connection>
<GID>72</GID>
<name>OUT_0</name></connection>
<intersection>-204 13</intersection>
<intersection>-180 7</intersection>
<intersection>-148 1</intersection>
<intersection>-114 3</intersection>
<intersection>-80 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121,-148,172.5,-148</points>
<connection>
<GID>124</GID>
<name>IN_1</name></connection>
<intersection>121 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>121,-114,172,-114</points>
<connection>
<GID>116</GID>
<name>IN_1</name></connection>
<intersection>121 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>121,-80,172,-80</points>
<connection>
<GID>91</GID>
<name>IN_1</name></connection>
<intersection>121 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>121,-180,173,-180</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<intersection>121 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>119,-204,121,-204</points>
<intersection>119 14</intersection>
<intersection>121 0</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>119,-277,119,-204</points>
<connection>
<GID>279</GID>
<name>IN_2</name></connection>
<intersection>-204 13</intersection></vsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124,-205,124,-68</points>
<connection>
<GID>73</GID>
<name>OUT_0</name></connection>
<intersection>-205 8</intersection>
<intersection>-183 7</intersection>
<intersection>-152 1</intersection>
<intersection>-118 3</intersection>
<intersection>-84 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>124,-152,172.5,-152</points>
<connection>
<GID>125</GID>
<name>IN_1</name></connection>
<intersection>124 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>124,-118,172,-118</points>
<connection>
<GID>117</GID>
<name>IN_1</name></connection>
<intersection>124 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>124,-84,172,-84</points>
<connection>
<GID>109</GID>
<name>IN_1</name></connection>
<intersection>124 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>124,-183,173,-183</points>
<connection>
<GID>133</GID>
<name>IN_0</name></connection>
<intersection>124 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>120,-205,124,-205</points>
<intersection>120 9</intersection>
<intersection>124 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>120,-277,120,-205</points>
<connection>
<GID>279</GID>
<name>IN_1</name></connection>
<intersection>-205 8</intersection></vsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>157,-205,157,-68</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>-205 5</intersection>
<intersection>-154 1</intersection>
<intersection>-120 2</intersection>
<intersection>-86 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>157,-154,172.5,-154</points>
<connection>
<GID>126</GID>
<name>IN_0</name></connection>
<intersection>157 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>157,-120,172,-120</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<intersection>157 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>157,-86,172,-86</points>
<connection>
<GID>110</GID>
<name>IN_0</name></connection>
<intersection>157 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>157,-205,178.5,-205</points>
<intersection>157 0</intersection>
<intersection>178.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>178.5,-239,178.5,-205</points>
<intersection>-239 7</intersection>
<intersection>-205 5</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>169.5,-239,178.5,-239</points>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<intersection>169.5 8</intersection>
<intersection>178.5 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>169.5,-239,169.5,-235</points>
<intersection>-239 7</intersection>
<intersection>-235 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>162.5,-235,169.5,-235</points>
<connection>
<GID>363</GID>
<name>IN_1</name></connection>
<intersection>169.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127,-206,127,-68</points>
<connection>
<GID>74</GID>
<name>OUT_0</name></connection>
<intersection>-206 8</intersection>
<intersection>-186 7</intersection>
<intersection>-156 1</intersection>
<intersection>-122 3</intersection>
<intersection>-88 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127,-156,172.5,-156</points>
<connection>
<GID>126</GID>
<name>IN_1</name></connection>
<intersection>127 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>127,-122,172,-122</points>
<connection>
<GID>118</GID>
<name>IN_1</name></connection>
<intersection>127 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>127,-88,172,-88</points>
<connection>
<GID>110</GID>
<name>IN_1</name></connection>
<intersection>127 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>127,-186,173,-186</points>
<connection>
<GID>134</GID>
<name>IN_0</name></connection>
<intersection>127 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>121,-206,127,-206</points>
<intersection>121 9</intersection>
<intersection>127 0</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>121,-277,121,-206</points>
<connection>
<GID>279</GID>
<name>IN_0</name></connection>
<intersection>-206 8</intersection></vsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>160,-204,160,-68</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<intersection>-204 5</intersection>
<intersection>-158 1</intersection>
<intersection>-124 2</intersection>
<intersection>-90 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>160,-158,172.5,-158</points>
<connection>
<GID>127</GID>
<name>IN_0</name></connection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>160,-124,172,-124</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>160,-90,172,-90</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<intersection>160 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>160,-204,181.5,-204</points>
<intersection>160 0</intersection>
<intersection>181.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>181.5,-247,181.5,-204</points>
<intersection>-247 7</intersection>
<intersection>-204 5</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>169.5,-247,181.5,-247</points>
<connection>
<GID>376</GID>
<name>IN_0</name></connection>
<intersection>169.5 8</intersection>
<intersection>181.5 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>169.5,-247,169.5,-243</points>
<intersection>-247 7</intersection>
<intersection>-243 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>162.5,-243,169.5,-243</points>
<connection>
<GID>349</GID>
<name>IN_1</name></connection>
<intersection>169.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130,-206,130,-68</points>
<connection>
<GID>75</GID>
<name>OUT_0</name></connection>
<intersection>-206 9</intersection>
<intersection>-189 7</intersection>
<intersection>-160 1</intersection>
<intersection>-126 3</intersection>
<intersection>-92 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>130,-160,172.5,-160</points>
<connection>
<GID>127</GID>
<name>IN_1</name></connection>
<intersection>130 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>130,-126,172,-126</points>
<connection>
<GID>119</GID>
<name>IN_1</name></connection>
<intersection>130 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>130,-92,172,-92</points>
<connection>
<GID>111</GID>
<name>IN_1</name></connection>
<intersection>130 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>130,-189,173,-189</points>
<connection>
<GID>135</GID>
<name>IN_0</name></connection>
<intersection>130 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>130,-206,136,-206</points>
<intersection>130 0</intersection>
<intersection>136 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>136,-277,136,-206</points>
<connection>
<GID>284</GID>
<name>IN_3</name></connection>
<intersection>-206 9</intersection></vsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163,-203,163,-68</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>-203 5</intersection>
<intersection>-162 1</intersection>
<intersection>-128 2</intersection>
<intersection>-94 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>163,-162,172.5,-162</points>
<connection>
<GID>128</GID>
<name>IN_0</name></connection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>163,-128,172,-128</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>163,-94,172,-94</points>
<connection>
<GID>112</GID>
<name>IN_0</name></connection>
<intersection>163 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>163,-203,184.5,-203</points>
<intersection>163 0</intersection>
<intersection>184.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>184.5,-255,184.5,-203</points>
<intersection>-255 7</intersection>
<intersection>-203 5</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>169.5,-255,184.5,-255</points>
<connection>
<GID>375</GID>
<name>IN_0</name></connection>
<intersection>169.5 8</intersection>
<intersection>184.5 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>169.5,-255,169.5,-251</points>
<intersection>-255 7</intersection>
<intersection>-251 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>162.5,-251,169.5,-251</points>
<connection>
<GID>351</GID>
<name>IN_1</name></connection>
<intersection>169.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,-205,133,-68</points>
<connection>
<GID>76</GID>
<name>OUT_0</name></connection>
<intersection>-205 9</intersection>
<intersection>-192 7</intersection>
<intersection>-164 1</intersection>
<intersection>-130 3</intersection>
<intersection>-96 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>133,-164,172.5,-164</points>
<connection>
<GID>128</GID>
<name>IN_1</name></connection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>133,-130,172,-130</points>
<connection>
<GID>120</GID>
<name>IN_1</name></connection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>133,-96,172,-96</points>
<connection>
<GID>112</GID>
<name>IN_1</name></connection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>133,-192,173,-192</points>
<connection>
<GID>136</GID>
<name>IN_0</name></connection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>133,-205,137,-205</points>
<intersection>133 0</intersection>
<intersection>137 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>137,-277,137,-205</points>
<connection>
<GID>284</GID>
<name>IN_2</name></connection>
<intersection>-205 9</intersection></vsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166,-202,166,-68</points>
<connection>
<GID>9</GID>
<name>OUT_0</name></connection>
<intersection>-202 5</intersection>
<intersection>-166 1</intersection>
<intersection>-132 2</intersection>
<intersection>-98 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>166,-166,172.5,-166</points>
<connection>
<GID>129</GID>
<name>IN_0</name></connection>
<intersection>166 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>166,-132,172,-132</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<intersection>166 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>166,-98,172,-98</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<intersection>166 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>166,-202,187.5,-202</points>
<intersection>166 0</intersection>
<intersection>187.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>187.5,-263,187.5,-202</points>
<intersection>-263 7</intersection>
<intersection>-202 5</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>169.5,-263,187.5,-263</points>
<connection>
<GID>374</GID>
<name>IN_0</name></connection>
<intersection>169.5 8</intersection>
<intersection>187.5 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>169.5,-263,169.5,-259</points>
<intersection>-263 7</intersection>
<intersection>-259 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>162.5,-259,169.5,-259</points>
<connection>
<GID>353</GID>
<name>IN_1</name></connection>
<intersection>169.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136,-204,136,-68</points>
<connection>
<GID>77</GID>
<name>OUT_0</name></connection>
<intersection>-204 9</intersection>
<intersection>-195 7</intersection>
<intersection>-168 1</intersection>
<intersection>-134 3</intersection>
<intersection>-100 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>136,-168,172.5,-168</points>
<connection>
<GID>129</GID>
<name>IN_1</name></connection>
<intersection>136 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>136,-134,172,-134</points>
<connection>
<GID>121</GID>
<name>IN_1</name></connection>
<intersection>136 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>136,-100,172,-100</points>
<connection>
<GID>113</GID>
<name>IN_1</name></connection>
<intersection>136 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>136,-195,173,-195</points>
<connection>
<GID>137</GID>
<name>IN_0</name></connection>
<intersection>136 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>136,-204,138,-204</points>
<intersection>136 0</intersection>
<intersection>138 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>138,-277,138,-204</points>
<connection>
<GID>284</GID>
<name>IN_1</name></connection>
<intersection>-204 9</intersection></vsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169,-201,169,-68</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>-201 4</intersection>
<intersection>-170 1</intersection>
<intersection>-136 2</intersection>
<intersection>-102 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>169,-170,172.5,-170</points>
<connection>
<GID>130</GID>
<name>IN_0</name></connection>
<intersection>169 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>169,-136,172,-136</points>
<connection>
<GID>122</GID>
<name>IN_0</name></connection>
<intersection>169 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>169,-102,172,-102</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>169 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>169,-201,190.5,-201</points>
<intersection>169 0</intersection>
<intersection>190.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>190.5,-271,190.5,-201</points>
<intersection>-271 7</intersection>
<intersection>-201 4</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>169.5,-271,190.5,-271</points>
<connection>
<GID>373</GID>
<name>IN_0</name></connection>
<intersection>169.5 8</intersection>
<intersection>190.5 6</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>169.5,-271,169.5,-267</points>
<intersection>-271 7</intersection>
<intersection>-267 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>162.5,-267,169.5,-267</points>
<connection>
<GID>355</GID>
<name>IN_1</name></connection>
<intersection>169.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139,-277,139,-68</points>
<connection>
<GID>78</GID>
<name>OUT_0</name></connection>
<connection>
<GID>284</GID>
<name>IN_0</name></connection>
<intersection>-198 5</intersection>
<intersection>-172 1</intersection>
<intersection>-138 2</intersection>
<intersection>-104 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>139,-172,172.5,-172</points>
<connection>
<GID>130</GID>
<name>IN_1</name></connection>
<intersection>139 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>139,-138,172,-138</points>
<connection>
<GID>122</GID>
<name>IN_1</name></connection>
<intersection>139 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>139,-104,172,-104</points>
<connection>
<GID>114</GID>
<name>IN_1</name></connection>
<intersection>139 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>139,-198,173,-198</points>
<connection>
<GID>140</GID>
<name>IN_0</name></connection>
<intersection>139 0</intersection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>131,-280,133,-280</points>
<connection>
<GID>284</GID>
<name>carry_out</name></connection>
<connection>
<GID>279</GID>
<name>carry_in</name></connection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155,-269,155,-268</points>
<intersection>-269 2</intersection>
<intersection>-268 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>155,-268,156.5,-268</points>
<connection>
<GID>355</GID>
<name>OUT</name></connection>
<intersection>155 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-269,155,-269</points>
<connection>
<GID>365</GID>
<name>IN_1</name></connection>
<intersection>155 0</intersection></hsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155,-272,155,-271</points>
<intersection>-272 2</intersection>
<intersection>-271 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>154,-271,155,-271</points>
<connection>
<GID>365</GID>
<name>IN_0</name></connection>
<intersection>155 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>155,-272,156.5,-272</points>
<connection>
<GID>356</GID>
<name>OUT</name></connection>
<intersection>155 0</intersection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155,-264,155,-263</points>
<intersection>-264 2</intersection>
<intersection>-263 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>154,-263,155,-263</points>
<connection>
<GID>366</GID>
<name>IN_0</name></connection>
<intersection>155 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>155,-264,156.5,-264</points>
<connection>
<GID>354</GID>
<name>OUT</name></connection>
<intersection>155 0</intersection></hsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155,-261,155,-260</points>
<intersection>-261 1</intersection>
<intersection>-260 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>154,-261,155,-261</points>
<connection>
<GID>366</GID>
<name>IN_1</name></connection>
<intersection>155 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>155,-260,156.5,-260</points>
<connection>
<GID>353</GID>
<name>OUT</name></connection>
<intersection>155 0</intersection></hsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155,-256,155,-255</points>
<intersection>-256 2</intersection>
<intersection>-255 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>154,-255,155,-255</points>
<connection>
<GID>367</GID>
<name>IN_0</name></connection>
<intersection>155 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>155,-256,156.5,-256</points>
<connection>
<GID>352</GID>
<name>OUT</name></connection>
<intersection>155 0</intersection></hsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155,-253,155,-252</points>
<intersection>-253 1</intersection>
<intersection>-252 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>154,-253,155,-253</points>
<connection>
<GID>367</GID>
<name>IN_1</name></connection>
<intersection>155 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>155,-252,156.5,-252</points>
<connection>
<GID>351</GID>
<name>OUT</name></connection>
<intersection>155 0</intersection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155,-248,155,-247</points>
<intersection>-248 2</intersection>
<intersection>-247 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>154,-247,155,-247</points>
<connection>
<GID>368</GID>
<name>IN_0</name></connection>
<intersection>155 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>155,-248,156.5,-248</points>
<connection>
<GID>350</GID>
<name>OUT</name></connection>
<intersection>155 0</intersection></hsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155,-245,155,-244</points>
<intersection>-245 1</intersection>
<intersection>-244 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>154,-245,155,-245</points>
<connection>
<GID>368</GID>
<name>IN_1</name></connection>
<intersection>155 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>155,-244,156.5,-244</points>
<connection>
<GID>349</GID>
<name>OUT</name></connection>
<intersection>155 0</intersection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155,-240,155,-239</points>
<intersection>-240 2</intersection>
<intersection>-239 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>154,-239,155,-239</points>
<connection>
<GID>369</GID>
<name>IN_0</name></connection>
<intersection>155 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>155,-240,156.5,-240</points>
<connection>
<GID>364</GID>
<name>OUT</name></connection>
<intersection>155 0</intersection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155,-237,155,-236</points>
<intersection>-237 1</intersection>
<intersection>-236 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>154,-237,155,-237</points>
<connection>
<GID>369</GID>
<name>IN_1</name></connection>
<intersection>155 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>155,-236,156.5,-236</points>
<connection>
<GID>363</GID>
<name>OUT</name></connection>
<intersection>155 0</intersection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155,-232,155,-231</points>
<intersection>-232 2</intersection>
<intersection>-231 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>154,-231,155,-231</points>
<connection>
<GID>370</GID>
<name>IN_0</name></connection>
<intersection>155 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>155,-232,156.5,-232</points>
<connection>
<GID>362</GID>
<name>OUT</name></connection>
<intersection>155 0</intersection></hsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155,-229,155,-228</points>
<intersection>-229 1</intersection>
<intersection>-228 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>154,-229,155,-229</points>
<connection>
<GID>370</GID>
<name>IN_1</name></connection>
<intersection>155 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>155,-228,156.5,-228</points>
<connection>
<GID>361</GID>
<name>OUT</name></connection>
<intersection>155 0</intersection></hsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155,-224,155,-223</points>
<intersection>-224 2</intersection>
<intersection>-223 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>154,-223,155,-223</points>
<connection>
<GID>371</GID>
<name>IN_0</name></connection>
<intersection>155 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>155,-224,156.5,-224</points>
<connection>
<GID>360</GID>
<name>OUT</name></connection>
<intersection>155 0</intersection></hsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155,-221,155,-220</points>
<intersection>-221 1</intersection>
<intersection>-220 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>154,-221,155,-221</points>
<connection>
<GID>371</GID>
<name>IN_1</name></connection>
<intersection>155 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>155,-220,156.5,-220</points>
<connection>
<GID>359</GID>
<name>OUT</name></connection>
<intersection>155 0</intersection></hsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155,-216,155,-215</points>
<intersection>-216 2</intersection>
<intersection>-215 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>154,-215,155,-215</points>
<connection>
<GID>372</GID>
<name>IN_0</name></connection>
<intersection>155 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>155,-216,156.5,-216</points>
<connection>
<GID>358</GID>
<name>OUT</name></connection>
<intersection>155 0</intersection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155,-213,155,-212</points>
<intersection>-213 1</intersection>
<intersection>-212 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>154,-213,155,-213</points>
<connection>
<GID>372</GID>
<name>IN_1</name></connection>
<intersection>155 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>155,-212,156.5,-212</points>
<connection>
<GID>357</GID>
<name>OUT</name></connection>
<intersection>155 0</intersection></hsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>146,-277,146,-270</points>
<connection>
<GID>284</GID>
<name>IN_B_0</name></connection>
<intersection>-270 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>146,-270,148,-270</points>
<connection>
<GID>365</GID>
<name>OUT</name></connection>
<intersection>146 0</intersection></hsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>162.5,-271,165.5,-271</points>
<connection>
<GID>356</GID>
<name>IN_1</name></connection>
<connection>
<GID>373</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>145,-277,145,-262</points>
<connection>
<GID>284</GID>
<name>IN_B_1</name></connection>
<intersection>-262 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>145,-262,148,-262</points>
<connection>
<GID>366</GID>
<name>OUT</name></connection>
<intersection>145 0</intersection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>162.5,-263,165.5,-263</points>
<connection>
<GID>354</GID>
<name>IN_1</name></connection>
<connection>
<GID>374</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>162.5,-255,165.5,-255</points>
<connection>
<GID>352</GID>
<name>IN_1</name></connection>
<connection>
<GID>375</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>162.5,-247,165.5,-247</points>
<connection>
<GID>350</GID>
<name>IN_1</name></connection>
<connection>
<GID>376</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>162.5,-231,165.5,-231</points>
<connection>
<GID>362</GID>
<name>IN_1</name></connection>
<connection>
<GID>164</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>162.5,-239,165.5,-239</points>
<connection>
<GID>364</GID>
<name>IN_1</name></connection>
<connection>
<GID>163</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>171</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>162.5,-223,165.5,-223</points>
<connection>
<GID>360</GID>
<name>IN_1</name></connection>
<connection>
<GID>165</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>162.5,-215,165.5,-215</points>
<connection>
<GID>358</GID>
<name>IN_1</name></connection>
<connection>
<GID>166</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>173</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144,-277,144,-254</points>
<connection>
<GID>284</GID>
<name>IN_B_2</name></connection>
<intersection>-254 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>144,-254,148,-254</points>
<connection>
<GID>367</GID>
<name>OUT</name></connection>
<intersection>144 0</intersection></hsegment></shape></wire>
<wire>
<ID>174</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>143,-277,143,-246</points>
<connection>
<GID>284</GID>
<name>IN_B_3</name></connection>
<intersection>-246 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>143,-246,148,-246</points>
<connection>
<GID>368</GID>
<name>OUT</name></connection>
<intersection>143 0</intersection></hsegment></shape></wire>
<wire>
<ID>175</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>128,-277,128,-238</points>
<connection>
<GID>279</GID>
<name>IN_B_0</name></connection>
<intersection>-238 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>128,-238,148,-238</points>
<connection>
<GID>369</GID>
<name>OUT</name></connection>
<intersection>128 0</intersection></hsegment></shape></wire>
<wire>
<ID>176</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127,-277,127,-230</points>
<connection>
<GID>279</GID>
<name>IN_B_1</name></connection>
<intersection>-230 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127,-230,148,-230</points>
<connection>
<GID>370</GID>
<name>OUT</name></connection>
<intersection>127 0</intersection></hsegment></shape></wire>
<wire>
<ID>177</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126,-277,126,-222</points>
<connection>
<GID>279</GID>
<name>IN_B_2</name></connection>
<intersection>-222 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>126,-222,148,-222</points>
<connection>
<GID>371</GID>
<name>OUT</name></connection>
<intersection>126 0</intersection></hsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,-277,125,-214</points>
<connection>
<GID>279</GID>
<name>IN_B_3</name></connection>
<intersection>-214 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>125,-214,148,-214</points>
<connection>
<GID>372</GID>
<name>OUT</name></connection>
<intersection>125 0</intersection></hsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>297,-120,297,-110</points>
<intersection>-120 1</intersection>
<intersection>-110 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>297,-120,298.5,-120</points>
<connection>
<GID>390</GID>
<name>N_in0</name></connection>
<intersection>297 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>288,-110,297,-110</points>
<connection>
<GID>381</GID>
<name>OUT</name></connection>
<intersection>297 0</intersection></hsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>295,-124,295,-117</points>
<intersection>-124 1</intersection>
<intersection>-117 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>295,-124,298.5,-124</points>
<connection>
<GID>391</GID>
<name>N_in0</name></connection>
<intersection>295 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>288,-117,295,-117</points>
<connection>
<GID>380</GID>
<name>OUT</name></connection>
<intersection>295 0</intersection></hsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>293,-128,293,-124</points>
<intersection>-128 1</intersection>
<intersection>-124 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>293,-128,298.5,-128</points>
<connection>
<GID>392</GID>
<name>N_in0</name></connection>
<intersection>293 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>288,-124,293,-124</points>
<connection>
<GID>379</GID>
<name>OUT</name></connection>
<intersection>293 0</intersection></hsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>293,-132,293,-131</points>
<intersection>-132 1</intersection>
<intersection>-131 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>293,-132,298.5,-132</points>
<connection>
<GID>393</GID>
<name>N_in0</name></connection>
<intersection>293 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>288,-131,293,-131</points>
<connection>
<GID>378</GID>
<name>OUT</name></connection>
<intersection>293 0</intersection></hsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>293,-137.5,293,-136</points>
<intersection>-137.5 2</intersection>
<intersection>-136 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>293,-136,298.5,-136</points>
<connection>
<GID>398</GID>
<name>N_in0</name></connection>
<intersection>293 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>288,-137.5,293,-137.5</points>
<connection>
<GID>385</GID>
<name>OUT</name></connection>
<intersection>293 0</intersection></hsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>293,-144.5,293,-140</points>
<intersection>-144.5 2</intersection>
<intersection>-140 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>293,-140,298.5,-140</points>
<connection>
<GID>399</GID>
<name>N_in0</name></connection>
<intersection>293 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>288,-144.5,293,-144.5</points>
<connection>
<GID>384</GID>
<name>OUT</name></connection>
<intersection>293 0</intersection></hsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>295,-151.5,295,-144</points>
<intersection>-151.5 2</intersection>
<intersection>-144 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>295,-144,298.5,-144</points>
<connection>
<GID>400</GID>
<name>N_in0</name></connection>
<intersection>295 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>288,-151.5,295,-151.5</points>
<connection>
<GID>383</GID>
<name>OUT</name></connection>
<intersection>295 0</intersection></hsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>297,-158.5,297,-148</points>
<intersection>-158.5 2</intersection>
<intersection>-148 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>297,-148,298.5,-148</points>
<connection>
<GID>401</GID>
<name>N_in0</name></connection>
<intersection>297 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>288,-158.5,297,-158.5</points>
<connection>
<GID>382</GID>
<name>OUT</name></connection>
<intersection>297 0</intersection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>0,235.418,1778,-681.582</PageViewport></page 3>
<page 4>
<PageViewport>0,235.418,1778,-681.582</PageViewport></page 4>
<page 5>
<PageViewport>0,235.418,1778,-681.582</PageViewport></page 5>
<page 6>
<PageViewport>0,235.418,1778,-681.582</PageViewport></page 6>
<page 7>
<PageViewport>0,235.418,1778,-681.582</PageViewport></page 7>
<page 8>
<PageViewport>0,235.418,1778,-681.582</PageViewport></page 8>
<page 9>
<PageViewport>0,235.418,1778,-681.582</PageViewport></page 9></circuit>